//: version "1.8.7"

module HalfAdd(B, A, S, C);
//: interface  /sz:(71, 88) /bd:[ Ti0>A(15/71) Ti1>B(54/71) Bo0<C(11/71) Bo1<S(58/71) ]
input B;    //: /sn:0 {0}(158,202)(250,202){1}
//: {2}(254,202)(323,202)(323,184)(331,184){3}
//: {4}(252,204)(252,248)(337,248){5}
input A;    //: /sn:0 {0}(157,155)(280,155){1}
//: {2}(284,155)(323,155)(323,179)(331,179){3}
//: {4}(282,157)(282,243)(337,243){5}
output C;    //: /sn:0 {0}(449,246)(358,246){1}
output S;    //: /sn:0 {0}(445,182)(352,182){1}
//: enddecls

  //: joint g4 (A) @(282, 155) /w:[ 2 -1 1 4 ]
  //: input g3 (B) @(156,202) /sn:0 /w:[ 0 ]
  //: input g2 (A) @(155,155) /sn:0 /w:[ 0 ]
  xor g1 (.I0(A), .I1(B), .Z(S));   //: @(342,182) /sn:0 /delay:" 2" /w:[ 3 3 1 ]
  //: output g6 (S) @(442,182) /sn:0 /w:[ 0 ]
  //: output g7 (C) @(446,246) /sn:0 /w:[ 0 ]
  //: joint g5 (B) @(252, 202) /w:[ 2 -1 1 4 ]
  and g0 (.I0(A), .I1(B), .Z(C));   //: @(348,246) /sn:0 /delay:" 1" /w:[ 5 5 1 ]

endmodule

module main;    //: root_module
wire [7:0] Z0;    //: /sn:0 {0}(488,272)(488,245)(488,245)(488,224){1}
wire [3:0] X0;    //: /sn:0 {0}(486,79)(486,131)(486,131)(486,141){1}
wire [3:0] Y0;    //: /sn:0 {0}(653,183)(574,183){1}
//: enddecls

  led g3 (.I(Z0));   //: @(488,279) /sn:0 /R:2 /w:[ 0 ] /type:3
  //: dip g2 (Y0) @(691,183) /sn:0 /R:3 /w:[ 0 ] /st:2
  //: dip g1 (X0) @(486,69) /sn:0 /w:[ 0 ] /st:5
  RCA g0 (.X(X0), .Y(Y0), .Z(Z0));   //: @(401, 142) /sz:(172, 81) /sn:0 /p:[ Ti0>1 Ri0>1 Bo0<1 ]

endmodule

module FullAdd(S, Cout, Cin, B, A);
//: interface  /sz:(83, 83) /bd:[ Ti0>A(19/83) Ti1>B(63/83) Ri0>Cin(42/83) Lo0<Cout(40/83) Bo0<S(43/83) ]
input B;    //: /sn:0 {0}(163,178)(214,178)(214,164)(224,164){1}
input A;    //: /sn:0 {0}(161,128)(224,128){1}
output Cout;    //: /sn:0 {0}(606,274)(567,274){1}
input Cin;    //: /sn:0 {0}(394,222)(182,222)(182,246)(165,246){1}
output S;    //: /sn:0 {0}(565,137)(500,137)(500,185)(484,185){1}
wire w3;    //: /sn:0 /dp:1 {0}(546,276)(318,276)(318,168)(308,168){1}
wire w2;    //: /sn:0 /dp:1 {0}(546,271)(494,271)(494,225)(484,225){1}
wire w5;    //: /sn:0 {0}(308,125)(386,125)(386,188)(394,188){1}
//: enddecls

  //: output g4 (S) @(562,137) /sn:0 /w:[ 0 ]
  //: output g3 (Cout) @(603,274) /sn:0 /w:[ 0 ]
  //: input g2 (Cin) @(163,246) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(161,178) /sn:0 /w:[ 0 ]
  HalfAdd g6 (.A(w5), .B(Cin), .S(S), .C(w2));   //: @(395, 174) /sz:(88, 62) /sn:0 /p:[ Li0>1 Li1>0 Ro0<1 Ro1<1 ]
  or g7 (.I0(w2), .I1(w3), .Z(Cout));   //: @(557,274) /sn:0 /w:[ 0 0 1 ]
  HalfAdd g5 (.A(A), .B(B), .S(w5), .C(w3));   //: @(225, 113) /sz:(82, 66) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<1 ]
  //: input g0 (A) @(159,128) /sn:0 /w:[ 0 ]

endmodule

module RCA(X, Z, Y);
//: interface  /sz:(172, 81) /bd:[ Ti0>X[3:0](89/180) Ri0>Y[3:0](41/81) Bo0<Z[7:0](92/180) ]
input [3:0] X;    //: /sn:0 {0}(163,26)(358,26){1}
//: {2}(359,26)(498,26){3}
//: {4}(499,26)(602,26){5}
//: {6}(603,26)(712,26){7}
//: {8}(713,26)(868,26){9}
output [7:0] Z;    //: /sn:0 {0}(925,791)(574,791)(574,826){1}
input [3:0] Y;    //: /sn:0 {0}(927,24)(927,58){1}
//: {2}(927,59)(927,111)(927,111)(927,140){3}
//: {4}(927,141)(927,243)(927,243)(927,359){5}
//: {6}(927,360)(927,545){7}
//: {8}(927,546)(927,622){9}
wire w32;    //: /sn:0 {0}(457,460)(416,460){1}
wire w6;    //: /sn:0 {0}(499,30)(499,74){1}
//: {2}(497,76)(429,76)(429,117){3}
//: {4}(427,119)(406,119)(406,347){5}
//: {6}(404,349)(386,349)(386,552){7}
//: {8}(406,351)(406,363){9}
//: {10}(429,121)(429,150){11}
//: {12}(499,78)(499,89)(499,89)(499,100){13}
wire B;    //: /sn:0 {0}(669,172)(669,226){1}
wire w7;    //: /sn:0 {0}(371,223)(371,127)(361,127)(361,117){1}
wire w46;    //: /sn:0 {0}(368,709)(368,867)(559,867)(559,832){1}
wire w16;    //: /sn:0 /dp:1 {0}(524,310)(524,342)(615,342)(615,413){1}
wire w14;    //: /sn:0 {0}(673,316)(673,340)(703,340)(703,858)(599,858)(599,832){1}
wire w19;    //: /sn:0 {0}(436,266)(483,266){1}
wire w15;    //: /sn:0 {0}(415,223)(415,194)(431,194)(431,171){1}
wire w4;    //: /sn:0 {0}(603,30)(603,74){1}
//: {2}(601,76)(580,76)(580,113){3}
//: {4}(578,115)(535,115)(535,347){5}
//: {6}(533,349)(511,349)(511,556){7}
//: {8}(535,351)(535,368){9}
//: {10}(580,117)(580,152){11}
//: {12}(603,78)(603,99){13}
wire w38;    //: /sn:0 {0}(409,667)(449,667){1}
wire A;    //: /sn:0 {0}(630,226)(630,168)(605,168)(605,120){1}
wire w0;    //: /sn:0 {0}(922,59)(720,59){1}
//: {2}(716,59)(610,59){3}
//: {4}(606,59)(506,59){5}
//: {6}(502,59)(364,59)(364,96){7}
//: {8}(504,61)(504,80)(504,80)(504,100){9}
//: {10}(608,61)(608,99){11}
//: {12}(718,61)(718,104){13}
wire w3;    //: /sn:0 {0}(922,141)(674,141){1}
//: {2}(670,141)(587,141){3}
//: {4}(583,141)(436,141){5}
//: {6}(432,141)(337,141)(337,152){7}
//: {8}(434,143)(434,150){9}
//: {10}(585,143)(585,152){11}
//: {12}(672,143)(672,151){13}
wire w43;    //: /sn:0 {0}(260,573)(260,622){1}
wire w21;    //: /sn:0 {0}(922,546)(647,546){1}
//: {2}(643,546)(518,546){3}
//: {4}(514,546)(393,546){5}
//: {6}(389,546)(263,546)(263,552){7}
//: {8}(391,548)(391,552){9}
//: {10}(516,548)(516,556){11}
//: {12}(645,548)(645,555){13}
wire w31;    //: /sn:0 {0}(344,624)(344,529)(243,529)(243,500){1}
wire w28;    //: /sn:0 {0}(642,576)(642,621){1}
wire w41;    //: /sn:0 {0}(534,669)(564,669)(564,723)(599,723)(599,711){1}
wire w36;    //: /sn:0 {0}(513,626)(513,577){1}
wire w23;    //: /sn:0 {0}(263,415)(263,394)(304,394)(304,384){1}
wire w24;    //: /sn:0 {0}(654,387)(654,413){1}
wire w20;    //: /sn:0 {0}(351,264)(328,264)(328,198)(238,198)(238,224){1}
wire w1;    //: /sn:0 {0}(713,30)(713,83){1}
//: {2}(711,85)(667,85)(667,117){3}
//: {4}(665,119)(652,119)(652,341){5}
//: {6}(650,343)(640,343)(640,555){7}
//: {8}(652,345)(652,366){9}
//: {10}(667,121)(667,151){11}
//: {12}(713,87)(713,104){13}
wire w25;    //: /sn:0 {0}(521,419)(521,396)(537,396)(537,389){1}
wire w35;    //: /sn:0 {0}(216,622)(216,589)(187,589)(187,456)(199,456){1}
wire w40;    //: /sn:0 {0}(388,573)(388,624){1}
wire w18;    //: /sn:0 {0}(477,419)(477,343)(395,343)(395,308){1}
wire w8;    //: /sn:0 {0}(359,30)(359,74){1}
//: {2}(357,76)(332,76)(332,114){3}
//: {4}(330,116)(302,116)(302,348){5}
//: {6}(300,350)(258,350)(258,552){7}
//: {8}(302,352)(302,363){9}
//: {10}(332,118)(332,152){11}
//: {12}(359,78)(359,96){13}
wire w30;    //: /sn:0 /dp:1 {0}(589,832)(589,870)(675,870)(675,536)(658,536)(658,503){1}
wire w22;    //: /sn:0 {0}(219,415)(219,363)(234,363)(234,314){1}
wire w17;    //: /sn:0 {0}(334,173)(334,176)(277,176)(277,224){1}
wire w44;    //: /sn:0 {0}(493,711)(493,878)(569,878)(569,832){1}
wire w11;    //: /sn:0 {0}(395,417)(395,393)(408,393)(408,384){1}
wire w12;    //: /sn:0 {0}(543,225)(543,189)(582,189)(582,173){1}
wire w2;    //: /sn:0 {0}(715,125)(715,131)(767,131)(767,849)(609,849)(609,832){1}
wire w10;    //: /sn:0 {0}(351,417)(351,340)(281,340)(281,314){1}
wire w27;    //: /sn:0 {0}(284,458)(338,458)(338,458)(331,458){1}
wire w13;    //: /sn:0 {0}(626,316)(626,332)(591,332)(591,268)(563,268){1}
wire w48;    //: /sn:0 {0}(240,707)(240,856)(549,856)(549,832){1}
wire w33;    //: /sn:0 {0}(469,626)(469,527)(375,527)(375,502){1}
wire w5;    //: /sn:0 {0}(501,225)(501,121){1}
wire w47;    //: /sn:0 {0}(196,663)(105,663)(105,846)(539,846)(539,832){1}
wire w29;    //: /sn:0 {0}(611,503)(611,519)(578,519)(578,462)(542,462){1}
wire w42;    //: /sn:0 {0}(281,665)(311,665)(311,665)(324,665){1}
wire w9;    //: /sn:0 {0}(922,360)(659,360){1}
//: {2}(655,360)(542,360){3}
//: {4}(538,360)(413,360){5}
//: {6}(409,360)(307,360)(307,363){7}
//: {8}(411,362)(411,363){9}
//: {10}(540,362)(540,368){11}
//: {12}(657,362)(657,366){13}
wire w39;    //: /sn:0 {0}(646,711)(646,880)(579,880)(579,832){1}
wire w26;    //: /sn:0 {0}(603,621)(603,534)(501,534)(501,504){1}
//: enddecls

  //: joint g61 (w8) @(302, 350) /w:[ -1 5 6 8 ]
  tran g4(.Z(w0), .I(Y[0]));   //: @(925,59) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:0
  //: joint g8 (w0) @(718, 59) /w:[ 1 -1 2 12 ]
  //: joint g58 (w21) @(516, 546) /w:[ 3 -1 4 10 ]
  and g55 (.I0(w21), .I1(w8), .Z(w43));   //: @(260,563) /sn:0 /R:3 /delay:" 1" /w:[ 7 7 0 ]
  tran g51(.Z(w21), .I(Y[3]));   //: @(925,546) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:0
  //: joint g37 (w9) @(657, 360) /w:[ 1 -1 2 12 ]
  tran g34(.Z(w9), .I(Y[2]));   //: @(925,360) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:0
  and g3 (.I0(w0), .I1(w1), .Z(w2));   //: @(715,115) /sn:0 /R:3 /delay:" 1" /w:[ 13 13 0 ]
  //: joint g13 (w0) @(504, 59) /w:[ 5 -1 6 8 ]
  FullAdd g65 (.B(w43), .A(w35), .Cin(w42), .Cout(w47), .S(w48));   //: @(197, 623) /sz:(83, 83) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>0 Lo0<0 Bo0<0 ]
  //: input g2 (X) @(161,26) /sn:0 /w:[ 0 ]
  //: joint g59 (w6) @(406, 349) /w:[ -1 5 6 8 ]
  concat g1 (.I0(w2), .I1(w14), .I2(w30), .I3(w39), .I4(w44), .I5(w46), .I6(w48), .I7(w47), .Z(Z));   //: @(574,827) /sn:0 /R:1 /w:[ 1 1 0 1 1 1 1 1 1 ] /dr:0
  FullAdd g64 (.B(w40), .A(w31), .Cin(w38), .Cout(w42), .S(w46));   //: @(325, 625) /sz:(83, 83) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  tran g11(.Z(w6), .I(X[2]));   //: @(499,24) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g16(.Z(w3), .I(Y[1]));   //: @(925,141) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:0
  and g50 (.I0(w21), .I1(w1), .Z(w28));   //: @(642,566) /sn:0 /R:3 /delay:" 1" /w:[ 13 7 0 ]
  //: joint g28 (w3) @(434, 141) /w:[ 5 -1 6 8 ]
  //: joint g10 (w0) @(608, 59) /w:[ 3 -1 4 10 ]
  //: output g19 (Z) @(922,791) /sn:0 /w:[ 0 ]
  and g27 (.I0(w3), .I1(w8), .Z(w17));   //: @(334,163) /sn:0 /R:3 /delay:" 1" /w:[ 7 11 0 ]
  //: joint g38 (w4) @(580, 115) /w:[ -1 3 4 10 ]
  and g6 (.I0(w0), .I1(w4), .Z(A));   //: @(605,110) /sn:0 /R:3 /delay:" 1" /w:[ 11 13 1 ]
  //: joint g57 (w4) @(535, 349) /w:[ -1 5 6 8 ]
  and g53 (.I0(w21), .I1(w4), .Z(w36));   //: @(513,567) /sn:0 /R:3 /delay:" 1" /w:[ 11 7 1 ]
  tran g7(.Z(w4), .I(X[1]));   //: @(603,24) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  and g9 (.I0(w0), .I1(w6), .Z(w5));   //: @(501,111) /sn:0 /R:3 /delay:" 1" /w:[ 9 13 1 ]
  HalfAdd g31 (.B(w17), .A(w20), .S(w10), .C(w22));   //: @(223, 225) /sz:(71, 88) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 Bo1<1 ]
  and g20 (.I0(w3), .I1(w4), .Z(w12));   //: @(582,163) /sn:0 /R:3 /delay:" 1" /w:[ 11 11 1 ]
  and g15 (.I0(w3), .I1(w1), .Z(B));   //: @(669,162) /sn:0 /R:3 /delay:" 1" /w:[ 13 11 0 ]
  and g39 (.I0(w9), .I1(w6), .Z(w11));   //: @(408,374) /sn:0 /R:3 /delay:" 1" /w:[ 9 9 1 ]
  FullAdd g48 (.B(w23), .A(w22), .Cin(w27), .Cout(w35), .S(w31));   //: @(200, 416) /sz:(83, 83) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<1 ]
  //: joint g43 (w9) @(411, 360) /w:[ 5 -1 6 8 ]
  HalfAdd g62 (.B(w28), .A(w26), .S(w39), .C(w41));   //: @(588, 622) /sz:(71, 88) /sn:0 /p:[ Ti0>1 Ti1>0 Bo0<0 Bo1<1 ]
  //: joint g29 (w8) @(359, 76) /w:[ -1 1 2 12 ]
  //: joint g25 (w3) @(585, 141) /w:[ 3 -1 4 10 ]
  //: joint g17 (w1) @(713, 85) /w:[ -1 1 2 12 ]
  FullAdd g63 (.B(w36), .A(w33), .Cin(w41), .Cout(w38), .S(w44));   //: @(450, 627) /sz:(83, 83) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g52 (w1) @(652, 343) /w:[ -1 5 6 8 ]
  and g42 (.I0(w9), .I1(w8), .Z(w23));   //: @(304,374) /sn:0 /R:3 /delay:" 1" /w:[ 7 9 1 ]
  //: joint g56 (w21) @(645, 546) /w:[ 1 -1 2 12 ]
  tran g5(.Z(w1), .I(X[0]));   //: @(713,24) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g14(.Z(w8), .I(X[3]));   //: @(359,24) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  FullAdd g47 (.B(w11), .A(w10), .Cin(w32), .Cout(w27), .S(w33));   //: @(332, 418) /sz:(83, 83) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<1 ]
  //: joint g44 (w8) @(332, 116) /w:[ -1 3 4 10 ]
  and g36 (.I0(w9), .I1(w4), .Z(w25));   //: @(537,379) /sn:0 /R:3 /delay:" 1" /w:[ 11 9 1 ]
  and g24 (.I0(w3), .I1(w6), .Z(w15));   //: @(431,161) /sn:0 /R:3 /delay:" 1" /w:[ 9 11 1 ]
  //: joint g21 (w4) @(603, 76) /w:[ -1 1 2 12 ]
  //: joint g41 (w6) @(429, 119) /w:[ -1 3 4 10 ]
  FullAdd g23 (.B(w12), .A(w5), .Cin(w13), .Cout(w19), .S(w16));   //: @(484, 226) /sz:(78, 83) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<0 ]
  //: joint g60 (w21) @(391, 546) /w:[ 5 -1 6 8 ]
  and g54 (.I0(w21), .I1(w6), .Z(w40));   //: @(388,563) /sn:0 /R:3 /delay:" 1" /w:[ 9 7 0 ]
  //: joint g40 (w9) @(540, 360) /w:[ 3 -1 4 10 ]
  HalfAdd g45 (.B(w24), .A(w16), .S(w30), .C(w29));   //: @(600, 414) /sz:(71, 88) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 Bo1<0 ]
  FullAdd g46 (.B(w25), .A(w18), .Cin(w29), .Cout(w32), .S(w26));   //: @(458, 420) /sz:(83, 83) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  //: joint g35 (w1) @(667, 119) /w:[ -1 3 4 10 ]
  //: joint g26 (w6) @(499, 76) /w:[ -1 1 2 12 ]
  //: joint g22 (w3) @(672, 141) /w:[ 1 -1 2 12 ]
  //: input g0 (Y) @(927,22) /sn:0 /R:3 /w:[ 0 ]
  and g12 (.I0(w0), .I1(w8), .Z(w7));   //: @(361,107) /sn:0 /R:3 /delay:" 1" /w:[ 7 13 1 ]
  HalfAdd g18 (.B(B), .A(A), .S(w14), .C(w13));   //: @(615, 227) /sz:(71, 88) /sn:0 /p:[ Ti0>1 Ti1>0 Bo0<0 Bo1<0 ]
  and g33 (.I0(w9), .I1(w1), .Z(w24));   //: @(654,377) /sn:0 /R:3 /delay:" 1" /w:[ 13 9 0 ]
  FullAdd g30 (.B(w15), .A(w7), .Cin(w19), .Cout(w20), .S(w18));   //: @(352, 224) /sz:(83, 83) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<1 ]

endmodule
