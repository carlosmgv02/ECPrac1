//: version "1.8.7"

module CPA4b(C0, C4, S, B, A);
//: interface  /sz:(104, 40) /bd:[ Ti0>B[3:0](67/104) Ti1>A[3:0](21/104) Ti2>A[3:0](21/104) Ti3>B[3:0](67/104) Ri0>C0(18/40) Ri1>C0(18/40) Lo0<C4(20/40) Lo1<C4(20/40) Bo0<S[3:0](46/104) Bo1<S[3:0](46/104) ]
input [3:0] B;    //: /sn:0 {0}(-59,44)(42,44){1}
//: {2}(43,44)(168,44){3}
//: {4}(169,44)(299,44){5}
//: {6}(300,44)(443,44){7}
//: {8}(444,44)(487,44){9}
input C0;    //: /sn:0 {0}(525,158)(465,158){1}
input [3:0] A;    //: /sn:0 {0}(-59,14)(-2,14){1}
//: {2}(-1,14)(124,14){3}
//: {4}(125,14)(255,14){5}
//: {6}(256,14)(399,14){7}
//: {8}(400,14)(495,14){9}
output C4;    //: /sn:0 {0}(-62,150)(-21,150){1}
output [3:0] S;    //: /sn:0 {0}(-115,321)(-23,321){1}
wire w6;    //: /sn:0 {0}(444,48)(444,115){1}
wire w7;    //: /sn:0 {0}(400,18)(400,115){1}
wire S1;    //: /sn:0 {0}(-17,316)(280,316)(280,198){1}
wire w16;    //: /sn:0 {0}(64,152)(105,152){1}
wire w4;    //: /sn:0 {0}(256,18)(256,113){1}
wire w0;    //: /sn:0 {0}(-1,18)(-1,109){1}
wire w3;    //: /sn:0 {0}(169,48)(169,111){1}
wire w23;    //: /sn:0 {0}(321,156)(380,156){1}
wire w24;    //: /sn:0 {0}(236,154)(190,154){1}
wire S0;    //: /sn:0 {0}(-17,306)(424,306)(424,200){1}
wire w8;    //: /sn:0 {0}(43,48)(43,109){1}
wire w2;    //: /sn:0 {0}(125,18)(125,111){1}
wire w5;    //: /sn:0 {0}(300,48)(300,113){1}
wire w9;    //: /sn:0 {0}(-17,336)(22,336)(22,194){1}
wire S2;    //: /sn:0 {0}(-17,326)(149,326)(149,196){1}
//: enddecls

  //: input g8 (C0) @(527,158) /sn:0 /R:2 /w:[ 0 ]
  tran g4(.Z(w3), .I(B[2]));   //: @(169,42) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: output g13 (C4) @(-59,150) /sn:0 /R:2 /w:[ 0 ]
  tran g3(.Z(w8), .I(B[3]));   //: @(43,42) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g2(.Z(w2), .I(A[2]));   //: @(125,12) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g1(.Z(w4), .I(A[1]));   //: @(256,12) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  FullAdd g28 (.B(w5), .A(w4), .Cin(w23), .Cout(w24), .S(S1));   //: @(237, 114) /sz:(83, 83) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<1 ]
  FullAdd g27 (.B(w3), .A(w2), .Cin(w24), .Cout(w16), .S(S2));   //: @(106, 112) /sz:(83, 83) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  tran g6(.Z(w7), .I(A[0]));   //: @(400,12) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g7(.Z(w6), .I(B[0]));   //: @(444,42) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: output g9 (S) @(-112,321) /sn:0 /R:2 /w:[ 0 ]
  //: input g15 (B) @(-61,44) /sn:0 /w:[ 0 ]
  FullAdd g29 (.B(w6), .A(w7), .Cin(C0), .Cout(w23), .S(S0));   //: @(381, 116) /sz:(83, 83) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  concat g17 (.I0(S0), .I1(S1), .I2(S2), .I3(w9), .Z(S));   //: @(-22,321) /sn:0 /R:2 /w:[ 0 0 0 0 1 ] /dr:0
  //: input g14 (A) @(-61,14) /sn:0 /w:[ 0 ]
  tran g5(.Z(w5), .I(B[1]));   //: @(300,42) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  FullAdd g26 (.B(w8), .A(w0), .Cin(w16), .Cout(C4), .S(w9));   //: @(-20, 110) /sz:(83, 83) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  tran g0(.Z(w0), .I(A[3]));   //: @(-1,12) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1

endmodule

module HalfAdd(B, A, S, C);
//: interface  /sz:(88, 71) /bd:[ Li0>A(16/71) Li1>B(55/71) Ro0<S(12/71) Ro1<C(59/71) ]
input B;    //: /sn:0 {0}(158,202)(250,202){1}
//: {2}(254,202)(320,202)(320,184)(328,184){3}
//: {4}(252,204)(252,248)(337,248){5}
input A;    //: /sn:0 {0}(157,155)(280,155){1}
//: {2}(284,155)(320,155)(320,179)(328,179){3}
//: {4}(282,157)(282,243)(337,243){5}
output C;    //: /sn:0 {0}(449,246)(358,246){1}
output S;    //: /sn:0 {0}(445,182)(349,182){1}
//: enddecls

  //: joint g4 (A) @(282, 155) /w:[ 2 -1 1 4 ]
  //: input g3 (B) @(156,202) /sn:0 /w:[ 0 ]
  //: input g2 (A) @(155,155) /sn:0 /w:[ 0 ]
  xor g1 (.I0(A), .I1(B), .Z(S));   //: @(339,182) /sn:0 /delay:" 2" /w:[ 3 3 1 ]
  //: output g6 (S) @(442,182) /sn:0 /w:[ 0 ]
  //: output g7 (C) @(446,246) /sn:0 /w:[ 0 ]
  //: joint g5 (B) @(252, 202) /w:[ 2 -1 1 4 ]
  and g0 (.I0(A), .I1(B), .Z(C));   //: @(348,246) /sn:0 /delay:" 1" /w:[ 5 5 1 ]

endmodule

module main;    //: root_module
wire [3:0] A0;    //: /sn:0 {0}(218,-11)(218,46)(218,46)(218,35){1}
wire w0;    //: /sn:0 {0}(372,79)(324,79)(324,79)(324,79){1}
wire [3:0] A;    //: /sn:0 /dp:1 {0}(54,-9)(54,35){1}
wire w1;    //: /sn:0 /dp:1 {0}(-31,77)(2,77)(2,77)(-4,77){1}
wire [3:0] w2;    //: /sn:0 /dp:1 {0}(150,146)(150,128)(150,128)(150,120){1}
//: enddecls

  led g4 (.I(w1));   //: @(-38,77) /sn:0 /R:1 /w:[ 0 ] /type:3
  //: switch g3 (w0) @(390,79) /sn:0 /R:2 /w:[ 0 ] /st:1
  //: dip g2 (A0) @(218,-21) /sn:0 /w:[ 0 ] /st:0
  //: dip g1 (A) @(54,-19) /sn:0 /w:[ 0 ] /st:9
  led g5 (.I(w2));   //: @(150,153) /sn:0 /R:2 /w:[ 0 ] /type:3
  CSA4b g0 (.B(A0), .A(A), .Cin(w0), .Cout(w1), .S(w2));   //: @(-3, 36) /sz:(326, 83) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]

endmodule

module FullAdd(S, Cout, Cin, B, A);
//: interface  /sz:(83, 83) /bd:[ Ti0>B(63/83) Ti1>A(19/83) Ti2>A(19/83) Ti3>B(63/83) Ri0>Cin(42/83) Ri1>Cin(42/83) Lo0<Cout(40/83) Lo1<Cout(40/83) Bo0<S(43/83) Bo1<S(43/83) ]
input B;    //: /sn:0 {0}(163,178)(214,178)(214,168)(224,168){1}
input A;    //: /sn:0 {0}(161,128)(192,128)(192,132)(224,132){1}
output Cout;    //: /sn:0 {0}(606,274)(567,274){1}
input Cin;    //: /sn:0 {0}(394,222)(182,222)(182,246)(165,246){1}
output S;    //: /sn:0 {0}(565,137)(500,137)(500,185)(484,185){1}
wire w3;    //: /sn:0 /dp:1 {0}(546,276)(318,276)(318,172)(308,172){1}
wire w2;    //: /sn:0 /dp:1 {0}(546,271)(494,271)(494,225)(484,225){1}
wire w5;    //: /sn:0 {0}(308,129)(386,129)(386,188)(394,188){1}
//: enddecls

  //: output g4 (S) @(562,137) /sn:0 /w:[ 0 ]
  //: output g3 (Cout) @(603,274) /sn:0 /w:[ 0 ]
  //: input g2 (Cin) @(163,246) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(161,178) /sn:0 /w:[ 0 ]
  HalfAdd g6 (.A(w5), .B(Cin), .S(S), .C(w2));   //: @(395, 174) /sz:(88, 62) /sn:0 /p:[ Li0>1 Li1>0 Ro0<1 Ro1<1 ]
  or g7 (.I0(w2), .I1(w3), .Z(Cout));   //: @(557,274) /sn:0 /delay:" 1" /w:[ 0 0 1 ]
  HalfAdd g5 (.A(A), .B(B), .S(w5), .C(w3));   //: @(225, 117) /sz:(82, 66) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<1 ]
  //: input g0 (A) @(159,128) /sn:0 /w:[ 0 ]

endmodule

module CSA4b(Cout, A, B, S, Cin);
//: interface  /sz:(326, 83) /bd:[ Ti0>A[3:0](57/326) Ti1>B[3:0](221/326) Ri0>Cin(43/83) Lo0<Cout(41/83) Bo0<S[3:0](153/326) ]
input [3:0] B;    //: /sn:0 {0}(176,96)(266,96)(266,96)(355,96){1}
//: {2}(356,96)(386,96)(386,96)(414,96){3}
//: {4}(415,96)(543,96){5}
supply0 w7;    //: /sn:0 {0}(555,164)(394,164){1}
supply1 w4;    //: /sn:0 {0}(559,225)(427,225)(427,246)(397,246){1}
input [3:0] A;    //: /sn:0 {0}(177,76)(262,76){1}
//: {2}(263,76)(287,76)(287,76)(309,76){3}
//: {4}(310,76)(535,76){5}
output Cout;    //: /sn:0 {0}(150,187)(181,187){1}
input Cin;    //: /sn:0 {0}(582,316)(504,316)(504,316)(457,316){1}
//: {2}(453,316)(380,316){3}
//: {4}(376,316)(305,316){5}
//: {6}(301,316)(210,316){7}
//: {8}(208,314)(208,238)(224,238)(224,128)(194,128)(194,164){9}
//: {10}(208,318)(208,344)(242,344){11}
//: {12}(303,318)(303,346)(320,346){13}
//: {14}(378,318)(378,346)(395,346){15}
//: {16}(455,318)(455,345)(471,345){17}
output [3:0] S;    //: /sn:0 {0}(582,403)(529,403){1}
wire [3:0] w6;    //: /sn:0 {0}(313,227)(313,193)(265,193){1}
//: {2}(263,191)(263,80){3}
//: {4}(261,193)(259,193){5}
wire [3:0] S1;    //: /sn:0 {0}(338,269)(338,275)(462,275){1}
//: {2}(463,275)(482,275){3}
//: {4}(483,275)(511,275){5}
//: {6}(512,275)(534,275){7}
//: {8}(535,275)(551,275){9}
wire w14;    //: /sn:0 {0}(265,357)(265,388)(523,388){1}
wire w19;    //: /sn:0 {0}(408,330)(408,314)(254,314)(254,276){1}
wire w15;    //: /sn:0 {0}(333,330)(333,319)(237,319)(237,276){1}
wire w3;    //: /sn:0 {0}(255,328)(255,323)(223,323)(223,276){1}
wire [3:0] w0;    //: /sn:0 {0}(356,145)(356,108)(356,108)(356,100){1}
wire S4;    //: /sn:0 {0}(353,330)(353,289)(483,289)(483,279){1}
wire w23;    //: /sn:0 {0}(484,329)(484,305)(269,305)(269,276){1}
wire [3:0] w1;    //: /sn:0 {0}(310,145)(310,88)(310,88)(310,80){1}
wire S0;    //: /sn:0 {0}(535,279)(535,296)(504,296)(504,329){1}
wire S5;    //: /sn:0 {0}(275,328)(275,284)(463,284)(463,279){1}
wire w18;    //: /sn:0 {0}(343,359)(343,398)(523,398){1}
wire w22;    //: /sn:0 {0}(418,359)(418,408)(523,408){1}
wire w11;    //: /sn:0 {0}(210,197)(272,197)(272,248)(291,248){1}
wire w10;    //: /sn:0 {0}(210,177)(278,177)(278,166)(288,166){1}
wire [3:0] w5;    //: /sn:0 {0}(359,227)(359,204)(415,204)(415,100){1}
wire S3;    //: /sn:0 {0}(428,330)(428,294)(512,294)(512,279){1}
wire [3:0] S2;    //: /sn:0 /dp:1 {0}(335,187)(335,217)(281,217)(281,272)(269,272){1}
//: {2}(268,272)(254,272){3}
//: {4}(253,272)(237,272){5}
//: {6}(236,272)(223,272){7}
//: {8}(222,272)(214,272){9}
wire w26;    //: /sn:0 {0}(494,358)(494,418)(523,418){1}
//: enddecls

  concat g8 (.I0(w26), .I1(w22), .I2(w18), .I3(w14), .Z(S));   //: @(528,403) /sn:0 /w:[ 1 1 1 1 1 ] /dr:0
  mux g4 (.I0(w3), .I1(S5), .S(Cin), .Z(w14));   //: @(265,344) /sn:0 /w:[ 0 0 11 0 ] /ss:136765592 /do:141333496
  //: output g3 (Cout) @(153,187) /sn:0 /R:2 /w:[ 0 ]
  //: input g13 (A) @(175,76) /sn:0 /w:[ 0 ]
  mux g2 (.I0(w10), .I1(w11), .S(Cin), .Z(Cout));   //: @(194,187) /sn:0 /R:3 /delay:" 1 1" /w:[ 0 0 9 1 ] /ss:-1514217216 /do:-1514217216
  CPA4b g1 (.A(w6), .B(w5), .C0(w4), .C4(w11), .S(S1));   //: @(292, 228) /sz:(104, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<0 ]
  //: input g16 (B) @(174,96) /sn:0 /w:[ 0 ]
  //: joint g11 (Cin) @(208, 316) /w:[ 7 8 -1 10 ]
  tran g28(.Z(S0), .I(S1[0]));   //: @(535,273) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: supply0 g10 (w7) @(561,164) /sn:0 /R:1 /w:[ 0 ]
  tran g32(.Z(S5), .I(S1[3]));   //: @(463,273) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g27(.Z(w23), .I(S2[0]));   //: @(269,270) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g19(.Z(w5), .I(B[3:0]));   //: @(415,94) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  mux g6 (.I0(w19), .I1(S3), .S(Cin), .Z(w22));   //: @(418,346) /sn:0 /w:[ 0 0 15 0 ] /ss:-1497440000 /do:-1497440000
  //: output g9 (S) @(579,403) /sn:0 /w:[ 0 ]
  mux g7 (.I0(w23), .I1(S0), .S(Cin), .Z(w26));   //: @(494,345) /sn:0 /w:[ 0 1 17 0 ] /ss:141689768 /do:141689744
  tran g31(.Z(S4), .I(S1[2]));   //: @(483,273) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g15(.Z(w6), .I(A[3:0]));   //: @(263,74) /sn:0 /R:1 /w:[ 3 1 2 ] /ss:1
  tran g20(.Z(w3), .I(S2[3]));   //: @(223,270) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  tran g25(.Z(w15), .I(S2[2]));   //: @(237,270) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  //: supply1 g29 (w4) @(559,236) /sn:0 /R:3 /w:[ 0 ]
  tran g17(.Z(w0), .I(B[3:0]));   //: @(356,94) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  mux g5 (.I0(w15), .I1(S4), .S(Cin), .Z(w18));   //: @(343,346) /sn:0 /w:[ 0 0 13 0 ] /ss:-1967136512 /do:-1933582080
  tran g14(.Z(w1), .I(A[3:0]));   //: @(310,74) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: input g21 (Cin) @(584,316) /sn:0 /R:2 /w:[ 0 ]
  //: joint g24 (Cin) @(303, 316) /w:[ 5 -1 6 12 ]
  //: joint g23 (Cin) @(378, 316) /w:[ 3 -1 4 14 ]
  tran g26(.Z(w19), .I(S2[1]));   //: @(254,270) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  CPA4b g0 (.A(w1), .B(w0), .C0(w7), .C4(w10), .S(S2));   //: @(289, 146) /sz:(104, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<0 ]
  //: joint g22 (Cin) @(455, 316) /w:[ 1 -1 2 16 ]
  //: joint g12 (w6) @(263, 193) /w:[ 1 2 4 -1 ]
  tran g30(.Z(S3), .I(S1[1]));   //: @(512,273) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1

endmodule
