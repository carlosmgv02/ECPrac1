//: version "1.8.7"

module PFA(A, Pi, Ci, S, Gi, B);
//: interface  /sz:(100, 97) /bd:[ Ti0>B(50/100) Ti1>A(14/100) Li0>Ci(46/97) Bo0<Gi(61/100) Ro0<Pi(67/97) Ro1<S(32/97) ]
input B;    //: /sn:0 {0}(184,223)(195,223){1}
//: {2}(199,223)(226,223)(226,207)(234,207){3}
//: {4}(197,225)(197,256){5}
//: {6}(199,258)(308,258){7}
//: {8}(197,260)(197,293)(309,293){9}
output Gi;    //: /sn:0 /dp:1 {0}(330,291)(354,291){1}
input A;    //: /sn:0 {0}(186,202)(214,202){1}
//: {2}(218,202)(234,202){3}
//: {4}(216,204)(216,251){5}
//: {6}(218,253)(308,253){7}
//: {8}(216,255)(216,288)(309,288){9}
output Pi;    //: /sn:0 /dp:1 {0}(329,256)(351,256){1}
input Ci;    //: /sn:0 /dp:1 {0}(305,227)(274,227)(274,241)(187,241){1}
output S;    //: /sn:0 {0}(358,225)(326,225){1}
wire w11;    //: /sn:0 {0}(255,205)(295,205)(295,222)(305,222){1}
//: enddecls

  //: input g4 (A) @(184,202) /sn:0 /w:[ 0 ]
  //: output g8 (Pi) @(348,256) /sn:0 /w:[ 1 ]
  xor g3 (.I0(A), .I1(B), .Z(w11));   //: @(245,205) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  xor g2 (.I0(w11), .I1(Ci), .Z(S));   //: @(316,225) /sn:0 /delay:" 2" /w:[ 1 0 1 ]
  or g1 (.I0(A), .I1(B), .Z(Pi));   //: @(319,256) /sn:0 /w:[ 7 7 0 ]
  //: joint g10 (A) @(216, 202) /w:[ 2 -1 1 4 ]
  //: input g6 (Ci) @(185,241) /sn:0 /w:[ 1 ]
  //: output g7 (S) @(355,225) /sn:0 /w:[ 0 ]
  //: output g9 (Gi) @(351,291) /sn:0 /w:[ 1 ]
  //: joint g12 (A) @(216, 253) /w:[ 6 5 -1 8 ]
  //: input g5 (B) @(182,223) /sn:0 /w:[ 0 ]
  //: joint g11 (B) @(197, 223) /w:[ 2 -1 1 4 ]
  and g0 (.I0(A), .I1(B), .Z(Gi));   //: @(320,291) /sn:0 /w:[ 9 9 0 ]
  //: joint g13 (B) @(197, 258) /w:[ 6 5 -1 8 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(202,175)(228,175)(228,200){1}
wire w7;    //: /sn:0 {0}(-28183,202)(-28183,212){1}
wire w4;    //: /sn:0 {0}(315,268)(345,268){1}
wire w3;    //: /sn:0 {0}(254,149)(264,149)(264,200){1}
wire w8;    //: /sn:0 {0}(181,247)(213,247){1}
wire w11;    //: /sn:0 {0}(275,321)(275,299){1}
wire w9;    //: /sn:0 {0}(345,233)(315,233){1}
//: enddecls

  led g4 (.I(w9));   //: @(352,233) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: switch g3 (w8) @(164,247) /sn:0 /w:[ 0 ] /st:1
  //: switch g2 (w7) @(-28183,189) /sn:0 /R:3 /w:[ 0 ] /st:0
  //: switch g1 (w6) @(185,175) /sn:0 /w:[ 0 ] /st:1
  led g6 (.I(w11));   //: @(275,328) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: switch g7 (w3) @(237,149) /sn:0 /w:[ 0 ] /st:0
  led g5 (.I(w4));   //: @(352,268) /sn:0 /R:3 /w:[ 1 ] /type:0
  PFA g0 (.B(w3), .A(w6), .Ci(w8), .Gi(w11), .Pi(w4), .S(w9));   //: @(214, 201) /sz:(100, 97) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Ro0<0 Ro1<1 ]

endmodule
