//: version "1.8.7"

module CLL(P1, G1, P0, G0, P3, C1, P2, C3, G2, C2, Cin, G3, C4);
//: interface  /sz:(383, 40) /bd:[ Ti0>G0(373/383) Ti1>P0(350/383) Ti2>G1(280/383) Ti3>P1(259/383) Ti4>G2(181/383) Ti5>P2(159/383) Ti6>G3(72/383) Ti7>P3(47/383) Ri0>Cin(22/40) To0<C1(294/383) To1<C2(199/383) To2<C3(96/383) Lo0<C4(21/40) ]
input G2;    //: /sn:0 {0}(82,119)(133,119){1}
//: {2}(137,119)(351,119)(351,90)(359,90){3}
//: {4}(135,117)(135,-32)(258,-32){5}
input P1;    //: /sn:0 {0}(95,192)(124,192){1}
//: {2}(128,192)(245,192)(245,186)(255,186){3}
//: {4}(126,190)(126,151){5}
//: {6}(128,149)(138,149)(138,150)(258,150){7}
//: {8}(126,147)(126,42){9}
//: {10}(128,40)(138,40)(138,41)(261,41){11}
//: {12}(126,38)(126,14){13}
output C3;    //: /sn:0 /dp:1 {0}(380,82)(410,82){1}
input G0;    //: /sn:0 /dp:1 {0}(354,256)(291,256)(291,273)(169,273){1}
//: {2}(167,271)(167,183){3}
//: {4}(169,181)(255,181){5}
//: {6}(167,179)(167,77){7}
//: {8}(169,75)(179,75)(179,76)(259,76){9}
//: {10}(167,73)(167,-101){11}
//: {12}(169,-103)(259,-103){13}
//: {14}(167,-105)(167,-144)(258,-144){15}
//: {16}(165,273)(100,273){17}
output C4;    //: /sn:0 {0}(423,-82)(383,-82){1}
output C2;    //: /sn:0 /dp:1 {0}(381,184)(419,184){1}
input Cin;    //: /sn:0 {0}(258,-149)(231,-149)(231,48){1}
//: {2}(233,50)(243,50)(243,51)(261,51){3}
//: {4}(231,52)(231,142){5}
//: {6}(233,144)(243,144)(243,145)(258,145){7}
//: {8}(231,146)(231,227){9}
//: {10}(233,229)(272,229){11}
//: {12}(231,231)(231,295)(92,295){13}
input P3;    //: /sn:0 {0}(258,-129)(78,-129)(78,-90){1}
//: {2}(80,-88)(259,-88){3}
//: {4}(78,-86)(78,-59){5}
//: {6}(80,-57)(259,-57){7}
//: {8}(78,-55)(78,-37){9}
//: {10}(80,-35)(250,-35)(250,-37)(258,-37){11}
//: {12}(76,-35)(65,-35){13}
input G1;    //: /sn:0 {0}(258,-139)(116,-139)(116,-100){1}
//: {2}(118,-98)(259,-98){3}
//: {4}(116,-96)(116,-69){5}
//: {6}(118,-67)(259,-67){7}
//: {8}(116,-65)(116,215){9}
//: {10}(118,217)(193,217){11}
//: {12}(197,217)(350,217)(350,189)(360,189){13}
//: {14}(195,215)(195,97)(260,97){15}
//: {16}(114,217)(96,217){17}
input G3;    //: /sn:0 {0}(66,-10)(352,-10)(352,-72)(362,-72){1}
output C1;    //: /sn:0 {0}(413,254)(375,254){1}
input P0;    //: /sn:0 {0}(261,46)(158,46)(158,45)(148,45){1}
//: {2}(146,43)(146,2){3}
//: {4}(146,47)(146,79){5}
//: {6}(148,81)(259,81){7}
//: {8}(146,83)(146,153){9}
//: {10}(148,155)(258,155){11}
//: {12}(146,157)(146,246){13}
//: {14}(148,248)(262,248)(262,234)(272,234){15}
//: {16}(144,248)(101,248){17}
input P2;    //: /sn:0 {0}(258,-134)(99,-134)(99,-95){1}
//: {2}(101,-93)(259,-93){3}
//: {4}(99,-91)(99,-64){5}
//: {6}(101,-62)(259,-62){7}
//: {8}(99,-60)(99,34){9}
//: {10}(101,36)(261,36){11}
//: {12}(99,38)(99,99){13}
//: {14}(101,101)(106,101){15}
//: {16}(110,101)(250,101)(250,102)(260,102){17}
//: {18}(108,99)(108,71)(259,71){19}
//: {20}(97,101)(80,101){21}
wire w6;    //: /sn:0 {0}(279,150)(355,150)(355,179)(360,179){1}
wire w13;    //: /sn:0 {0}(279,-34)(345,-34)(345,-77)(362,-77){1}
wire w7;    //: /sn:0 /dp:1 {0}(362,-87)(305,-87)(305,-96)(280,-96){1}
wire w4;    //: /sn:0 {0}(293,232)(344,232)(344,251)(354,251){1}
wire w3;    //: /sn:0 {0}(359,85)(342,85)(342,100)(281,100){1}
wire w0;    //: /sn:0 /dp:1 {0}(359,75)(337,75)(337,43)(282,43){1}
wire w10;    //: /sn:0 {0}(279,-139)(311,-139)(311,-92)(362,-92){1}
wire w1;    //: /sn:0 /dp:1 {0}(359,80)(325,80)(325,76)(280,76){1}
wire w11;    //: /sn:0 {0}(280,-62)(341,-62)(341,-82)(362,-82){1}
wire w5;    //: /sn:0 {0}(276,184)(360,184){1}
//: enddecls

  and g8 (.I0(Cin), .I1(P0), .Z(w4));   //: @(283,232) /sn:0 /w:[ 11 15 0 ]
  //: input g4 (P1) @(93,192) /sn:0 /w:[ 0 ]
  //: joint g44 (G1) @(116, 217) /w:[ 10 9 16 -1 ]
  and g16 (.I0(Cin), .I1(P1), .I2(P0), .Z(w6));   //: @(269,150) /sn:0 /w:[ 7 7 11 0 ]
  //: input g3 (G1) @(94,217) /sn:0 /w:[ 17 ]
  //: joint g47 (P2) @(99, -62) /w:[ 6 5 -1 8 ]
  //: joint g26 (P2) @(108, 101) /w:[ 16 18 15 -1 ]
  //: joint g17 (Cin) @(231, 144) /w:[ 6 5 -1 8 ]
  //: input g2 (P0) @(99,248) /sn:0 /w:[ 17 ]
  //: joint g30 (Cin) @(231, 50) /w:[ 2 1 -1 4 ]
  and g23 (.I0(G1), .I1(P2), .Z(w3));   //: @(271,100) /sn:0 /w:[ 15 17 1 ]
  //: joint g24 (G1) @(195, 217) /w:[ 12 14 11 -1 ]
  //: input g1 (G0) @(98,273) /sn:0 /w:[ 17 ]
  //: input g39 (P3) @(63,-35) /sn:0 /w:[ 13 ]
  and g29 (.I0(P2), .I1(P1), .I2(P0), .I3(Cin), .Z(w0));   //: @(272,43) /sn:0 /w:[ 11 11 0 3 1 ]
  //: joint g51 (P2) @(99, -93) /w:[ 2 1 -1 4 ]
  //: joint g18 (P1) @(126, 192) /w:[ 2 4 1 -1 ]
  and g25 (.I0(P2), .I1(G0), .I2(P0), .Z(w1));   //: @(270,76) /sn:0 /w:[ 19 9 7 1 ]
  //: output g10 (C1) @(410,254) /sn:0 /w:[ 0 ]
  and g49 (.I0(Cin), .I1(G0), .I2(G1), .I3(P2), .I4(P3), .Z(w10));   //: @(269,-139) /sn:0 /w:[ 0 15 0 0 0 0 ]
  //: input g6 (P2) @(78,101) /sn:0 /w:[ 21 ]
  //: joint g50 (P3) @(78, -88) /w:[ 2 1 -1 4 ]
  //: output g35 (C3) @(407,82) /sn:0 /w:[ 1 ]
  //: joint g9 (Cin) @(231, 229) /w:[ 10 9 -1 12 ]
  or g7 (.I0(w4), .I1(G0), .Z(C1));   //: @(365,254) /sn:0 /w:[ 1 0 1 ]
  //: joint g31 (P0) @(146, 45) /w:[ 1 2 -1 4 ]
  or g22 (.I0(w0), .I1(w1), .I2(w3), .I3(G2), .Z(C3));   //: @(370,82) /sn:0 /w:[ 0 0 0 3 0 ]
  //: joint g33 (P2) @(99, 101) /w:[ 14 13 20 -1 ]
  or g36 (.I0(w10), .I1(w7), .I2(w11), .I3(w13), .I4(G3), .Z(C4));   //: @(373,-82) /sn:0 /w:[ 1 0 1 1 1 1 ]
  //: joint g41 (G2) @(135, 119) /w:[ 2 4 1 -1 ]
  and g45 (.I0(G0), .I1(G1), .I2(P2), .I3(P3), .Z(w7));   //: @(270,-96) /sn:0 /w:[ 13 3 3 3 1 ]
  and g40 (.I0(P3), .I1(G2), .Z(w13));   //: @(269,-34) /sn:0 /w:[ 11 5 0 ]
  and g42 (.I0(G1), .I1(P2), .I2(P3), .Z(w11));   //: @(270,-62) /sn:0 /w:[ 7 7 7 0 ]
  //: joint g52 (G1) @(116, -98) /w:[ 2 1 -1 4 ]
  and g12 (.I0(G0), .I1(P1), .Z(w5));   //: @(266,184) /sn:0 /w:[ 5 3 0 ]
  //: joint g34 (P2) @(99, 36) /w:[ 10 9 -1 12 ]
  //: joint g28 (P0) @(146, 81) /w:[ 6 5 -1 8 ]
  //: joint g46 (P3) @(78, -57) /w:[ 6 5 -1 8 ]
  //: joint g14 (G0) @(167, 181) /w:[ 4 6 -1 3 ]
  or g11 (.I0(w6), .I1(w5), .I2(G1), .Z(C2));   //: @(371,184) /sn:0 /w:[ 1 1 13 0 ]
  //: input g5 (G2) @(80,119) /sn:0 /w:[ 0 ]
  //: output g21 (C2) @(416,184) /sn:0 /w:[ 1 ]
  //: joint g19 (P1) @(126, 149) /w:[ 6 8 -1 5 ]
  //: joint g32 (P1) @(126, 40) /w:[ 10 12 -1 9 ]
  //: joint g20 (P0) @(146, 155) /w:[ 10 9 -1 12 ]
  //: joint g15 (P0) @(146, 248) /w:[ 14 13 16 -1 ]
  //: input g0 (Cin) @(90,295) /sn:0 /w:[ 13 ]
  //: input g38 (G3) @(64,-10) /sn:0 /w:[ 0 ]
  //: joint g43 (P3) @(78, -35) /w:[ 10 9 12 -1 ]
  //: joint g27 (G0) @(167, 75) /w:[ 8 10 -1 7 ]
  //: joint g48 (G1) @(116, -67) /w:[ 6 5 -1 8 ]
  //: output g37 (C4) @(420,-82) /sn:0 /w:[ 0 ]
  //: joint g13 (G0) @(167, 273) /w:[ 1 2 16 -1 ]
  //: joint g53 (G0) @(167, -103) /w:[ 12 14 -1 11 ]

endmodule

module PFA(Pi, S, Ci, B, Gi, A);
//: interface  /sz:(40, 40) /bd:[ Li0>A(8/40) Li1>B(23/40) Li2>Ci(37/40) Ro0<S(12/40) Ro1<Pi(26/40) Ro2<Gi(37/40) ]
input B;    //: /sn:0 {0}(206,145)(223,145){1}
//: {2}(227,145)(269,145)(269,133)(279,133){3}
//: {4}(225,147)(225,188){5}
//: {6}(227,190)(354,190){7}
//: {8}(225,192)(225,229)(356,229){9}
output Gi;    //: /sn:0 {0}(435,225)(387,225)(387,227)(377,227){1}
input A;    //: /sn:0 {0}(205,117)(246,117){1}
//: {2}(250,117)(269,117)(269,128)(279,128){3}
//: {4}(248,119)(248,183){5}
//: {6}(250,185)(354,185){7}
//: {8}(248,187)(248,224)(356,224){9}
output Pi;    //: /sn:0 /dp:1 {0}(375,188)(422,188)(422,187)(432,187){1}
input Ci;    //: /sn:0 /dp:1 {0}(351,146)(314,146)(314,174)(204,174){1}
output S;    //: /sn:0 /dp:1 {0}(372,144)(423,144)(423,145)(433,145){1}
wire w2;    //: /sn:0 {0}(300,131)(341,131)(341,141)(351,141){1}
//: enddecls

  or g8 (.I0(A), .I1(B), .Z(Pi));   //: @(365,188) /sn:0 /w:[ 7 7 0 ]
  //: output g4 (Pi) @(429,187) /sn:0 /w:[ 1 ]
  //: output g3 (S) @(430,145) /sn:0 /w:[ 1 ]
  //: input g2 (Ci) @(202,174) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(204,145) /sn:0 /w:[ 0 ]
  //: joint g10 (A) @(248, 117) /w:[ 2 -1 1 4 ]
  xor g6 (.I0(A), .I1(B), .Z(w2));   //: @(290,131) /sn:0 /w:[ 3 3 0 ]
  and g9 (.I0(A), .I1(B), .Z(Gi));   //: @(367,227) /sn:0 /w:[ 9 9 1 ]
  xor g7 (.I0(w2), .I1(Ci), .Z(S));   //: @(362,144) /sn:0 /w:[ 1 0 0 ]
  //: joint g12 (B) @(225, 145) /w:[ 2 -1 1 4 ]
  //: joint g11 (A) @(248, 185) /w:[ 6 5 -1 8 ]
  //: output g5 (Gi) @(432,225) /sn:0 /w:[ 0 ]
  //: input g0 (A) @(203,117) /sn:0 /w:[ 0 ]
  //: joint g13 (B) @(225, 190) /w:[ 6 5 -1 8 ]

endmodule

module main;    //: root_module
wire [3:0] w4;    //: /sn:0 {0}(323,232)(323,222){1}
wire [3:0] w3;    //: /sn:0 {0}(285,232)(285,222){1}
wire [3:0] w0;    //: /sn:0 {0}(285,114)(285,124){1}
wire [3:0] w1;    //: /sn:0 {0}(322,114)(322,124){1}
wire w2;    //: /sn:0 {0}(434,159)(424,159){1}
wire [3:0] w5;    //: /sn:0 {0}(374,232)(374,222){1}
//: enddecls

  CLA g0 (.B(w1), .A(w0), .Cin(w2), .P(w5), .G(w4), .S(w3));   //: @(261, 125) /sz:(162, 96) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Bo0<1 Bo1<1 Bo2<1 ]

endmodule

module CLA(A, B, Cin);
//: interface  /sz:(162, 96) /bd:[ Ti0>A[3:0](24/162) Ti1>B[3:0](61/162) Ri0>Cin(34/96) Bo0<S[3:0](24/162) Bo1<G[3:0](62/162) Bo2<P[3:0](113/162) ]
input [3:0] B;    //: /sn:0 {0}(117,75)(205,75){1}
//: {2}(206,75)(306,75){3}
//: {4}(307,75)(406,75){5}
//: {6}(407,75)(498,75){7}
//: {8}(499,75)(558,75){9}
input [3:0] A;    //: /sn:0 {0}(126,58)(175,58){1}
//: {2}(176,58)(277,58){3}
//: {4}(278,58)(378,58){5}
//: {6}(379,58)(469,58){7}
//: {8}(470,58)(557,58){9}
input Cin;    //: /sn:0 {0}(574,109)(557,109){1}
//: {2}(553,109)(526,109)(526,120){3}
//: {4}(555,111)(555,238)(538,238){5}
wire w16;    //: /sn:0 {0}(412,164)(412,205)(413,205)(413,215){1}
wire w13;    //: /sn:0 {0}(407,122)(407,79){1}
wire w6;    //: /sn:0 {0}(278,123)(278,62){1}
wire w7;    //: /sn:0 {0}(307,123)(307,79){1}
wire w4;    //: /sn:0 {0}(201,164)(201,215){1}
wire w22;    //: /sn:0 {0}(505,165)(505,205)(504,205)(504,215){1}
wire w3;    //: /sn:0 {0}(174,164)(174,174){1}
wire w0;    //: /sn:0 {0}(176,122)(176,62){1}
wire w20;    //: /sn:0 /dp:1 {0}(448,215)(448,112)(433,112)(433,122){1}
wire w19;    //: /sn:0 {0}(499,120)(499,79){1}
wire w18;    //: /sn:0 {0}(470,120)(470,62){1}
wire w12;    //: /sn:0 {0}(379,122)(379,62){1}
wire w23;    //: /sn:0 {0}(526,165)(526,205)(527,205)(527,215){1}
wire w10;    //: /sn:0 {0}(313,165)(313,215){1}
wire w21;    //: /sn:0 {0}(478,165)(478,175){1}
wire w1;    //: /sn:0 {0}(206,122)(206,79){1}
wire w8;    //: /sn:0 /dp:1 {0}(250,215)(250,112)(234,112)(234,122){1}
wire w17;    //: /sn:0 {0}(433,164)(433,205)(434,205)(434,215){1}
wire w14;    //: /sn:0 /dp:1 {0}(353,215)(353,113)(334,113)(334,123){1}
wire w2;    //: /sn:0 {0}(143,237)(153,237){1}
wire w11;    //: /sn:0 {0}(334,165)(334,205)(335,205)(335,215){1}
wire w15;    //: /sn:0 {0}(386,164)(386,174){1}
wire w5;    //: /sn:0 {0}(225,164)(225,205)(226,205)(226,215){1}
wire w9;    //: /sn:0 {0}(286,165)(286,175){1}
//: enddecls

  tran g8(.Z(w0), .I(A[3]));   //: @(176,56) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: input g4 (A) @(559,58) /sn:0 /R:2 /w:[ 9 ]
  CLL g16 (.P3(w4), .G3(w5), .P2(w10), .G2(w11), .P1(w16), .G1(w17), .P0(w22), .G0(w23), .Cin(Cin), .C3(w8), .C2(w14), .C1(w20), .C4(w2));   //: @(154, 216) /sz:(383, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>5 To0<0 To1<0 To2<0 Lo0<1 ]
  PFA g3 (.Ci(Cin), .B(w19), .A(w18), .G0(w23), .P0(w22), .S(w21));   //: @(455, 121) /sz:(77, 43) /sn:0 /p:[ Ti0>3 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  PFA g2 (.Ci(w20), .B(w13), .A(w12), .G1(w17), .P1(w16), .S(w15));   //: @(364, 123) /sz:(75, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  PFA g1 (.Ci(w14), .B(w7), .A(w6), .G2(w11), .P2(w10), .S(w9));   //: @(263, 124) /sz:(77, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  tran g10(.Z(w19), .I(B[0]));   //: @(499,73) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g6(.Z(w12), .I(A[1]));   //: @(379,56) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g9 (B) @(560,75) /sn:0 /R:2 /w:[ 9 ]
  tran g7(.Z(w6), .I(A[2]));   //: @(278,56) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g12(.Z(w7), .I(B[2]));   //: @(307,73) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: input g14 (Cin) @(576,109) /sn:0 /R:2 /w:[ 0 ]
  tran g11(.Z(w13), .I(B[1]));   //: @(407,73) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g5(.Z(w18), .I(A[0]));   //: @(470,56) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: joint g15 (Cin) @(555, 109) /w:[ 1 -1 2 4 ]
  PFA g0 (.Ci(w8), .B(w1), .A(w0), .G3(w5), .P3(w4), .S(w3));   //: @(160, 123) /sz:(80, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  tran g13(.Z(w1), .I(B[3]));   //: @(206,73) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1

endmodule
