//: version "1.8.7"

module PFA2();
//: interface  /sz:(40, 40) /bd:[ ]
wire w6;    //: /sn:0 {0}(203,112)(223,112)(223,112)(247,112){1}
//: {2}(249,110)(249,100)(298,100)(298,90)(327,90){3}
//: {4}(249,114)(249,172)(353,172){5}
wire w7;    //: /sn:0 {0}(203,151)(375,151)(375,119)(402,119){1}
wire w0;    //: /sn:0 {0}(499,59)(472,59)(472,88)(377,88){1}
//: {2}(373,88)(348,88){3}
//: {4}(375,90)(375,114)(402,114){5}
wire w8;    //: /sn:0 {0}(499,170)(374,170){1}
wire w2;    //: /sn:0 {0}(499,117)(423,117){1}
wire w5;    //: /sn:0 {0}(203,70)(274,70){1}
//: {2}(278,70)(298,70)(298,85)(327,85){3}
//: {4}(276,72)(276,167)(353,167){5}
//: enddecls

  xor g4 (.I0(w0), .I1(w7), .Z(w2));   //: @(413,117) /sn:0 /delay:" 2" /w:[ 5 1 1 ]
  //: switch g8 (w7) @(186,151) /sn:0 /w:[ 0 ] /st:0
  xor g3 (.I0(w5), .I1(w6), .Z(w0));   //: @(338,88) /sn:0 /delay:" 2" /w:[ 3 3 3 ]
  //: joint g2 (w0) @(375, 88) /w:[ 1 -1 2 4 ]
  //: joint g1 (w6) @(249, 112) /w:[ -1 2 1 4 ]
  led g11 (.I(w8));   //: @(506,170) /sn:0 /R:3 /w:[ 0 ] /type:3
  led g10 (.I(w2));   //: @(506,117) /sn:0 /R:3 /w:[ 0 ] /type:3
  //: switch g6 (w5) @(186,70) /sn:0 /w:[ 0 ] /st:0
  //: switch g7 (w6) @(186,112) /sn:0 /w:[ 0 ] /st:0
  led g9 (.I(w0));   //: @(506,59) /sn:0 /R:3 /w:[ 0 ] /type:3
  and g5 (.I0(w5), .I1(w6), .Z(w8));   //: @(364,170) /sn:0 /delay:" 1" /w:[ 5 5 1 ]
  //: joint g0 (w5) @(276, 70) /w:[ 2 -1 1 4 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(137,102)(157,102)(157,102)(181,102){1}
//: {2}(183,100)(183,90)(232,90)(232,80)(261,80){3}
//: {4}(183,104)(183,167)(286,167){5}
wire w7;    //: /sn:0 {0}(137,141)(309,141)(309,109)(336,109){1}
wire w0;    //: /sn:0 {0}(433,49)(406,49)(406,78)(311,78){1}
//: {2}(307,78)(282,78){3}
//: {4}(309,80)(309,104)(336,104){5}
wire w8;    //: /sn:0 {0}(433,160)(369,160)(369,165)(307,165){1}
wire w2;    //: /sn:0 {0}(433,107)(357,107){1}
wire w5;    //: /sn:0 {0}(137,60)(208,60){1}
//: {2}(212,60)(232,60)(232,75)(261,75){3}
//: {4}(210,62)(210,162)(286,162){5}
//: enddecls

  xor g4 (.I0(w0), .I1(w7), .Z(w2));   //: @(347,107) /sn:0 /delay:" 2" /w:[ 5 1 1 ]
  //: switch g8 (w7) @(120,141) /sn:0 /w:[ 0 ] /st:1
  xor g3 (.I0(w5), .I1(w6), .Z(w0));   //: @(272,78) /sn:0 /delay:" 2" /w:[ 3 3 3 ]
  //: joint g2 (w0) @(309, 78) /w:[ 1 -1 2 4 ]
  //: joint g1 (w6) @(183, 102) /w:[ -1 2 1 4 ]
  led g11 (.I(w8));   //: @(440,160) /sn:0 /R:3 /w:[ 0 ] /type:3
  led g10 (.I(w2));   //: @(440,107) /sn:0 /R:3 /w:[ 0 ] /type:3
  //: switch g6 (w5) @(120,60) /sn:0 /w:[ 0 ] /st:0
  //: switch g7 (w6) @(120,102) /sn:0 /w:[ 0 ] /st:1
  led g9 (.I(w0));   //: @(440,49) /sn:0 /R:3 /w:[ 0 ] /type:3
  and g5 (.I0(w5), .I1(w6), .Z(w8));   //: @(297,165) /sn:0 /delay:" 1" /w:[ 5 5 1 ]
  //: joint g0 (w5) @(210, 60) /w:[ 2 -1 1 4 ]

endmodule
