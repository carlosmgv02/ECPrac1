//: version "1.8.7"

module CLL(P1, G1, P0, G0, P3, C1, P2, C3, GG, G2, C2, Cin, G3, C4, PG);
//: interface  /sz:(385, 86) /bd:[ Ti0>G0(374/385) Ti1>P0(351/385) Ti2>G1(281/385) Ti3>P1(260/385) Ti4>G2(181/385) Ti5>P2(159/385) Ti6>G3(72/385) Ti7>P3(47/385) Ri0>Cin(47/86) To0<C1(295/385) To1<C2(200/385) To2<C3(96/385) Lo0<C4(45/86) Bo0<GG(331/385) Bo1<PG(271/385) ]
input G2;    //: {0}(82,119)(133,119){1}
//: {2}(137,119)(317,119){3}
//: {4}(321,119)(351,119)(351,90)(359,90){5}
//: {6}(319,117)(319,-1)(367,-1){7}
//: {8}(135,117)(135,-32)(258,-32){9}
output GG;    //: /sn:0 {0}(595,3)(585,3)(585,18)(667,18)(667,26)(652,-7)(569,-7){1}
input P1;    //: /sn:0 {0}(-47,-29)(-30,-29)(-30,10)(7,10)(7,155){1}
//: {2}(9,157)(101,157)(101,190){3}
//: {4}(103,192)(124,192){5}
//: {6}(128,192)(205,192){7}
//: {8}(209,192)(245,192)(245,186)(255,186){9}
//: {10}(207,190)(207,-51)(496,-51){11}
//: {12}(126,190)(126,151){13}
//: {14}(128,149)(138,149)(138,150)(258,150){15}
//: {16}(126,147)(126,42){17}
//: {18}(128,40)(138,40)(138,41)(261,41){19}
//: {20}(126,38)(126,14){21}
//: {22}(99,192)(95,192){23}
//: {24}(5,157)(-5,157){25}
output C3;    //: /sn:0 /dp:1 {0}(380,82)(410,82){1}
output PG;    //: /sn:0 /dp:1 {0}(-68,-31)(-82,-31)(-82,94)(-101,94){1}
input G0;    //: /sn:0 /dp:1 {0}(499,278)(456,278){1}
//: {2}(454,276)(454,-56)(496,-56){3}
//: {4}(452,278)(436,278)(436,273)(169,273){5}
//: {6}(167,271)(167,183){7}
//: {8}(169,181)(255,181){9}
//: {10}(167,179)(167,77){11}
//: {12}(169,75)(179,75)(179,76)(259,76){13}
//: {14}(167,73)(167,-101){15}
//: {16}(169,-103)(259,-103){17}
//: {18}(167,-105)(167,-144)(258,-144){19}
//: {20}(165,273)(100,273){21}
output C4;    //: /sn:0 {0}(423,-82)(383,-82){1}
output C2;    //: /sn:0 /dp:1 {0}(381,184)(419,184){1}
input Cin;    //: /sn:0 {0}(258,-149)(231,-149)(231,48){1}
//: {2}(233,50)(243,50)(243,51)(261,51){3}
//: {4}(231,52)(231,142){5}
//: {6}(233,144)(243,144)(243,145)(258,145){7}
//: {8}(231,146)(231,227){9}
//: {10}(233,229)(272,229){11}
//: {12}(231,231)(231,295)(92,295){13}
input P3;    //: /sn:0 {0}(390,28)(378,28)(378,19)(354,19)(354,-4){1}
//: {2}(356,-6)(367,-6){3}
//: {4}(352,-6)(335,-6){5}
//: {6}(333,-8)(333,-29)(432,-29)(432,-46)(496,-46){7}
//: {8}(331,-6)(237,-6)(237,-33){9}
//: {10}(239,-35)(250,-35)(250,-37)(258,-37){11}
//: {12}(235,-35)(80,-35){13}
//: {14}(78,-37)(78,-55){15}
//: {16}(80,-57)(259,-57){17}
//: {18}(78,-59)(78,-86){19}
//: {20}(80,-88)(259,-88){21}
//: {22}(78,-90)(78,-129)(258,-129){23}
//: {24}(76,-35)(44,-35)(44,-44){25}
//: {26}(44,-48)(44,-57)(39,-57){27}
//: {28}(42,-46)(-2,-46)(-2,-39)(-47,-39){29}
input G1;    //: /sn:0 {0}(390,38)(299,38)(299,215){1}
//: {2}(301,217)(350,217)(350,189)(360,189){3}
//: {4}(297,217)(197,217){5}
//: {6}(195,215)(195,97)(260,97){7}
//: {8}(193,217)(118,217){9}
//: {10}(116,215)(116,-65){11}
//: {12}(118,-67)(259,-67){13}
//: {14}(116,-69)(116,-96){15}
//: {16}(118,-98)(259,-98){17}
//: {18}(116,-100)(116,-139)(258,-139){19}
//: {20}(114,217)(96,217){21}
input G3;    //: /sn:0 {0}(548,-14)(483,-14)(483,-17)(320,-17){1}
//: {2}(318,-19)(318,-72)(362,-72){3}
//: {4}(316,-17)(306,-17)(306,-16)(27,-16){5}
input P0;    //: /sn:0 {0}(-47,-24)(-17,-24)(-17,29)(-11,29)(-11,219){1}
//: {2}(-9,221)(115,221)(115,246){3}
//: {4}(117,248)(144,248){5}
//: {6}(148,248)(262,248)(262,234)(272,234){7}
//: {8}(146,246)(146,157){9}
//: {10}(148,155)(258,155){11}
//: {12}(146,153)(146,83){13}
//: {14}(148,81)(259,81){15}
//: {16}(146,79)(146,47){17}
//: {18}(148,45)(158,45)(158,46)(261,46){19}
//: {20}(146,43)(146,2){21}
//: {22}(113,248)(101,248){23}
//: {24}(-13,221)(-26,221){25}
output C1;    //: /sn:0 {0}(657,257)(652,257)(652,276)(520,276){1}
input P2;    //: /sn:0 {0}(-47,-34)(-1,-34)(-1,1)(87,1)(87,99){1}
//: {2}(89,101)(97,101){3}
//: {4}(101,101)(106,101){5}
//: {6}(110,101)(177,101){7}
//: {8}(181,101)(244,101){9}
//: {10}(248,101)(250,101)(250,102)(260,102){11}
//: {12}(246,99)(246,33)(390,33){13}
//: {14}(179,99)(179,-23)(470,-23)(470,-41)(496,-41){15}
//: {16}(108,99)(108,71)(259,71){17}
//: {18}(99,99)(99,38){19}
//: {20}(101,36)(261,36){21}
//: {22}(99,34)(99,-60){23}
//: {24}(101,-62)(259,-62){25}
//: {26}(99,-64)(99,-91){27}
//: {28}(101,-93)(259,-93){29}
//: {30}(99,-95)(99,-134)(258,-134){31}
//: {32}(85,101)(80,101){33}
wire w16;    //: /sn:0 {0}(517,-49)(538,-49)(538,1)(548,1){1}
wire w6;    //: /sn:0 {0}(279,150)(355,150)(355,179)(360,179){1}
wire w13;    //: /sn:0 {0}(279,-34)(345,-34)(345,-77)(362,-77){1}
wire w7;    //: /sn:0 /dp:1 {0}(362,-87)(305,-87)(305,-96)(280,-96){1}
wire w4;    //: /sn:0 {0}(293,232)(489,232)(489,273)(499,273){1}
wire w3;    //: /sn:0 {0}(359,85)(342,85)(342,100)(281,100){1}
wire w0;    //: /sn:0 /dp:1 {0}(359,75)(337,75)(337,43)(282,43){1}
wire w12;    //: /sn:0 {0}(548,-4)(501,-4)(501,33)(411,33){1}
wire w10;    //: /sn:0 {0}(279,-139)(311,-139)(311,-92)(362,-92){1}
wire w1;    //: /sn:0 /dp:1 {0}(359,80)(325,80)(325,76)(280,76){1}
wire w11;    //: /sn:0 {0}(280,-62)(341,-62)(341,-82)(362,-82){1}
wire w15;    //: /sn:0 {0}(388,-3)(489,-3)(489,-9)(548,-9){1}
wire w5;    //: /sn:0 {0}(276,184)(360,184){1}
//: enddecls

  //: joint g75 (G0) @(454, 278) /w:[ 1 2 4 -1 ]
  and g8 (.I0(Cin), .I1(P0), .Z(w4));   //: @(283,232) /sn:0 /delay:" 3" /w:[ 11 7 0 ]
  //: input g4 (P1) @(93,192) /sn:0 /w:[ 23 ]
  //: joint g44 (G1) @(116, 217) /w:[ 9 10 20 -1 ]
  and g16 (.I0(Cin), .I1(P1), .I2(P0), .Z(w6));   //: @(269,150) /sn:0 /delay:" 3" /w:[ 7 15 11 0 ]
  //: input g3 (G1) @(94,217) /sn:0 /w:[ 21 ]
  //: joint g47 (P2) @(99, -62) /w:[ 24 26 -1 23 ]
  //: joint g26 (P2) @(108, 101) /w:[ 6 16 5 -1 ]
  //: joint g17 (Cin) @(231, 144) /w:[ 6 5 -1 8 ]
  //: input g2 (P0) @(99,248) /sn:0 /w:[ 23 ]
  //: joint g74 (P1) @(207, 192) /w:[ 8 10 7 -1 ]
  //: joint g30 (Cin) @(231, 50) /w:[ 2 1 -1 4 ]
  and g23 (.I0(G1), .I1(P2), .Z(w3));   //: @(271,100) /sn:0 /delay:" 3" /w:[ 7 11 1 ]
  //: joint g24 (G1) @(195, 217) /w:[ 5 6 8 -1 ]
  //: input g1 (G0) @(98,273) /sn:0 /w:[ 21 ]
  //: input g39 (P3) @(37,-57) /sn:0 /w:[ 27 ]
  //: joint g60 (P0) @(115, 248) /w:[ 4 3 22 -1 ]
  and g29 (.I0(P2), .I1(P1), .I2(P0), .I3(Cin), .Z(w0));   //: @(272,43) /sn:0 /delay:" 3" /w:[ 21 19 19 3 1 ]
  //: joint g51 (P2) @(99, -93) /w:[ 28 30 -1 27 ]
  //: joint g70 (G1) @(299, 217) /w:[ 2 1 4 -1 ]
  //: joint g18 (P1) @(126, 192) /w:[ 6 12 5 -1 ]
  //: joint g65 (P3) @(237, -35) /w:[ 10 -1 12 9 ]
  and g25 (.I0(P2), .I1(G0), .I2(P0), .Z(w1));   //: @(270,76) /sn:0 /delay:" 3" /w:[ 17 13 15 1 ]
  //: output g10 (C1) @(654,257) /sn:0 /w:[ 0 ]
  or g64 (.I0(G3), .I1(w15), .I2(w12), .I3(w16), .Z(GG));   //: @(559,-7) /sn:0 /delay:" 3" /w:[ 0 1 0 1 1 ]
  //: joint g72 (P3) @(333, -6) /w:[ 5 6 8 -1 ]
  and g49 (.I0(Cin), .I1(G0), .I2(G1), .I3(P2), .I4(P3), .Z(w10));   //: @(269,-139) /sn:0 /delay:" 3" /w:[ 0 19 19 31 23 0 ]
  //: input g6 (P2) @(78,101) /sn:0 /w:[ 33 ]
  //: joint g50 (P3) @(78, -88) /w:[ 20 22 -1 19 ]
  //: joint g73 (P2) @(179, 101) /w:[ 8 14 7 -1 ]
  //: joint g68 (P3) @(354, -6) /w:[ 2 -1 4 1 ]
  //: joint g58 (P1) @(101, 192) /w:[ 4 3 22 -1 ]
  //: joint g56 (P3) @(44, -46) /w:[ -1 26 28 25 ]
  //: output g35 (C3) @(407,82) /sn:0 /w:[ 1 ]
  //: joint g9 (Cin) @(231, 229) /w:[ 10 9 -1 12 ]
  or g7 (.I0(w4), .I1(G0), .Z(C1));   //: @(510,276) /sn:0 /delay:" 3" /w:[ 1 0 1 ]
  and g71 (.I0(P3), .I1(P2), .I2(G1), .Z(w12));   //: @(401,33) /sn:0 /delay:" 3" /w:[ 0 13 0 1 ]
  //: joint g59 (P1) @(7, 157) /w:[ 2 1 24 -1 ]
  //: joint g31 (P0) @(146, 45) /w:[ 18 20 -1 17 ]
  or g22 (.I0(w0), .I1(w1), .I2(w3), .I3(G2), .Z(C3));   //: @(370,82) /sn:0 /delay:" 3" /w:[ 0 0 0 5 0 ]
  and g67 (.I0(P3), .I1(G2), .Z(w15));   //: @(378,-3) /sn:0 /delay:" 3" /w:[ 3 7 0 ]
  //: output g54 (GG) @(592,3) /sn:0 /w:[ 0 ]
  //: joint g33 (P2) @(99, 101) /w:[ 4 18 3 -1 ]
  or g36 (.I0(w10), .I1(w7), .I2(w11), .I3(w13), .I4(G3), .Z(C4));   //: @(373,-82) /sn:0 /delay:" 3" /w:[ 1 0 1 1 3 1 ]
  //: joint g41 (G2) @(135, 119) /w:[ 2 8 1 -1 ]
  and g45 (.I0(G0), .I1(G1), .I2(P2), .I3(P3), .Z(w7));   //: @(270,-96) /sn:0 /delay:" 3" /w:[ 17 17 29 21 1 ]
  //: joint g69 (P2) @(246, 101) /w:[ 10 12 9 -1 ]
  and g40 (.I0(P3), .I1(G2), .Z(w13));   //: @(269,-34) /sn:0 /delay:" 3" /w:[ 11 9 0 ]
  and g42 (.I0(G1), .I1(P2), .I2(P3), .Z(w11));   //: @(270,-62) /sn:0 /delay:" 3" /w:[ 13 25 17 0 ]
  //: joint g52 (G1) @(116, -98) /w:[ 16 18 -1 15 ]
  //: joint g66 (G2) @(319, 119) /w:[ 4 6 3 -1 ]
  and g12 (.I0(G0), .I1(P1), .Z(w5));   //: @(266,184) /sn:0 /delay:" 3" /w:[ 9 9 0 ]
  //: joint g57 (P2) @(87, 101) /w:[ 2 1 32 -1 ]
  //: joint g34 (P2) @(99, 36) /w:[ 20 22 -1 19 ]
  //: joint g28 (P0) @(146, 81) /w:[ 14 16 -1 13 ]
  //: joint g46 (P3) @(78, -57) /w:[ 16 18 -1 15 ]
  //: joint g14 (G0) @(167, 181) /w:[ 8 10 -1 7 ]
  or g11 (.I0(w6), .I1(w5), .I2(G1), .Z(C2));   //: @(371,184) /sn:0 /delay:" 3" /w:[ 1 1 3 0 ]
  //: input g5 (G2) @(80,119) /sn:0 /w:[ 0 ]
  //: joint g61 (P0) @(-11, 221) /w:[ 2 1 24 -1 ]
  //: output g21 (C2) @(416,184) /sn:0 /w:[ 1 ]
  //: joint g19 (P1) @(126, 149) /w:[ 14 16 -1 13 ]
  //: joint g32 (P1) @(126, 40) /w:[ 18 20 -1 17 ]
  //: joint g20 (P0) @(146, 155) /w:[ 10 12 -1 9 ]
  //: joint g63 (G3) @(318, -17) /w:[ 1 2 4 -1 ]
  //: joint g15 (P0) @(146, 248) /w:[ 6 8 5 -1 ]
  //: input g0 (Cin) @(90,295) /sn:0 /w:[ 13 ]
  //: input g38 (G3) @(25,-16) /sn:0 /w:[ 5 ]
  //: joint g43 (P3) @(78, -35) /w:[ 13 14 24 -1 ]
  //: joint g27 (G0) @(167, 75) /w:[ 12 14 -1 11 ]
  //: joint g48 (G1) @(116, -67) /w:[ 12 14 -1 11 ]
  and g62 (.I0(P0), .I1(P1), .I2(P2), .I3(P3), .Z(PG));   //: @(-58,-31) /sn:0 /R:2 /delay:" 3" /w:[ 0 0 0 29 0 ]
  //: output g37 (C4) @(420,-82) /sn:0 /w:[ 0 ]
  //: output g55 (PG) @(-98,94) /sn:0 /R:2 /w:[ 1 ]
  and g76 (.I0(G0), .I1(P1), .I2(P3), .I3(P2), .Z(w16));   //: @(507,-49) /sn:0 /delay:" 3" /w:[ 3 11 7 15 0 ]
  //: joint g13 (G0) @(167, 273) /w:[ 5 6 20 -1 ]
  //: joint g53 (G0) @(167, -103) /w:[ 16 18 -1 15 ]

endmodule

module PFA(Pi, S, Ci, B, Gi, A);
//: interface  /sz:(40, 40) /bd:[ Li0>A(8/40) Li1>B(23/40) Li2>Ci(37/40) Ro0<S(12/40) Ro1<Pi(26/40) Ro2<Gi(37/40) ]
input B;    //: /sn:0 {0}(206,145)(223,145){1}
//: {2}(227,145)(269,145)(269,133)(279,133){3}
//: {4}(225,147)(225,188){5}
//: {6}(227,190)(354,190){7}
//: {8}(225,192)(225,229)(356,229){9}
output Gi;    //: /sn:0 {0}(435,225)(387,225)(387,227)(377,227){1}
input A;    //: /sn:0 {0}(205,117)(246,117){1}
//: {2}(250,117)(269,117)(269,128)(279,128){3}
//: {4}(248,119)(248,183){5}
//: {6}(250,185)(354,185){7}
//: {8}(248,187)(248,224)(356,224){9}
output Pi;    //: /sn:0 /dp:1 {0}(375,188)(422,188)(422,187)(432,187){1}
input Ci;    //: /sn:0 /dp:1 {0}(352,146)(315,146)(315,174)(204,174){1}
output S;    //: /sn:0 /dp:1 {0}(373,144)(424,144)(424,145)(433,145){1}
wire w2;    //: /sn:0 {0}(300,131)(342,131)(342,141)(352,141){1}
//: enddecls

  or g8 (.I0(A), .I1(B), .Z(Pi));   //: @(365,188) /sn:0 /delay:" 3" /w:[ 7 7 0 ]
  //: output g4 (Pi) @(429,187) /sn:0 /w:[ 1 ]
  //: output g3 (S) @(430,145) /sn:0 /w:[ 1 ]
  //: input g2 (Ci) @(202,174) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(204,145) /sn:0 /w:[ 0 ]
  //: joint g10 (A) @(248, 117) /w:[ 2 -1 1 4 ]
  xor g6 (.I0(A), .I1(B), .Z(w2));   //: @(290,131) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  and g9 (.I0(A), .I1(B), .Z(Gi));   //: @(367,227) /sn:0 /delay:" 3" /w:[ 9 9 1 ]
  xor g7 (.I0(w2), .I1(Ci), .Z(S));   //: @(363,144) /sn:0 /delay:" 4" /w:[ 1 0 0 ]
  //: joint g12 (B) @(225, 145) /w:[ 2 -1 1 4 ]
  //: joint g11 (A) @(248, 185) /w:[ 6 5 -1 8 ]
  //: output g5 (Gi) @(432,225) /sn:0 /w:[ 0 ]
  //: input g0 (A) @(203,117) /sn:0 /w:[ 0 ]
  //: joint g13 (B) @(225, 190) /w:[ 6 5 -1 8 ]

endmodule

module main;    //: root_module
wire w16;    //: /sn:0 {0}(252,267)(252,238)(176,238){1}
//: {2}(174,236)(174,185)(180,185){3}
//: {4}(174,240)(174,245){5}
wire w6;    //: /sn:0 /dp:1 {0}(283,-71)(283,-25)(497,-25)(497,140)(472,140){1}
wire w7;    //: /sn:0 /dp:1 {0}(273,-71)(273,22)(349,22)(349,127)(366,127)(366,142)(356,142){1}
wire w34;    //: /sn:0 {0}(472,181)(483,181)(483,195)(426,195)(426,267){1}
wire w4;    //: /sn:0 {0}(135,168)(158,168)(158,229)(99,229)(99,267){1}
wire w0;    //: /sn:0 {0}(61,187)(54,187)(54,204)(148,204)(148,267){1}
wire w3;    //: /sn:0 {0}(135,187)(146,187)(146,201)(124,201)(124,267){1}
wire w22;    //: /sn:0 {0}(246,185)(257,185)(257,199)(233,199)(233,267){1}
wire w20;    //: /sn:0 {0}(180,163)(158,163)(158,76){1}
wire w29;    //: /sn:0 {0}(356,164)(376,164)(376,221)(312,221)(312,267){1}
wire [3:0] w37;    //: /sn:0 {0}(-105,72)(-105,102)(28,102){1}
//: {2}(29,102)(166,102){3}
//: {4}(167,102)(276,102){5}
//: {6}(277,102)(383,102){7}
//: {8}(384,102)(531,102){9}
wire w12;    //: /sn:0 {0}(387,416)(387,365)(383,365)(383,355){1}
wire w18;    //: /sn:0 {0}(51,313)(-23,313)(-23,281){1}
wire w10;    //: /sn:0 {0}(263,-71)(263,17)(236,17)(236,130)(256,130)(256,145)(246,145){1}
wire w21;    //: /sn:0 {0}(180,139)(167,139)(167,106){1}
wire w1;    //: /sn:0 {0}(61,163)(-9,163)(-9,76){1}
wire w32;    //: /sn:0 {0}(401,158)(376,158)(376,76){1}
wire w8;    //: /sn:0 {0}(211,267)(211,213)(266,213){1}
//: {2}(268,211)(268,167)(246,167){3}
//: {4}(268,215)(268,227){5}
wire w17;    //: /sn:0 {0}(347,267)(347,229)(283,229)(283,182)(292,182){1}
wire w27;    //: /sn:0 {0}(292,135)(277,135)(277,106){1}
wire w28;    //: /sn:0 {0}(356,182)(367,182)(367,196)(333,196)(333,267){1}
wire w33;    //: /sn:0 {0}(401,134)(384,134)(384,106){1}
wire w35;    //: /sn:0 {0}(472,163)(498,163)(498,242){1}
//: {2}(496,244)(414,244)(414,243)(404,243){3}
//: {4}(402,241)(402,236){5}
//: {6}(402,245)(402,256)(403,256)(403,267){7}
//: {8}(498,246)(498,254){9}
wire w14;    //: /sn:0 {0}(438,315)(530,315)(530,215){1}
//: {2}(532,213)(579,213)(579,252){3}
//: {4}(528,213)(390,213)(390,181)(401,181){5}
wire w2;    //: /sn:0 {0}(61,139)(29,139)(29,106){1}
wire [3:0] w11;    //: /sn:0 /dp:1 {0}(383,-84)(268,-84)(268,-77){1}
wire w5;    //: /sn:0 {0}(135,145)(141,145)(141,-25)(253,-25)(253,-71){1}
wire [3:0] w38;    //: /sn:0 {0}(568,72)(376,72){1}
//: {2}(375,72)(265,72){3}
//: {4}(264,72)(158,72){5}
//: {6}(157,72)(-9,72){7}
//: {8}(-10,72)(-44,72)(-44,38){9}
wire w9;    //: /sn:0 {0}(240,420)(323,420)(323,355){1}
wire w26;    //: /sn:0 {0}(292,159)(265,159)(265,76){1}
//: enddecls

  PFA g4 (.A(w33), .B(w32), .Ci(w14), .S(w6), .Pi(w35), .Gi(w34));   //: @(402, 121) /sz:(69, 65) /sn:0 /p:[ Li0>0 Li1>0 Li2>5 Ro0<1 Ro1<0 Ro2<0 ]
  tran g8(.Z(w27), .I(w37[1]));   //: @(277,100) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  PFA g3 (.A(w27), .B(w26), .Ci(w17), .S(w7), .Pi(w29), .Gi(w28));   //: @(293, 123) /sz:(62, 64) /sn:0 /p:[ Li0>0 Li1>0 Li2>1 Ro0<1 Ro1<0 Ro2<0 ]
  //: joint g16 (w35) @(498, 244) /w:[ -1 1 2 8 ]
  //: joint g17 (w35) @(402, 243) /w:[ 3 4 -1 6 ]
  PFA g2 (.A(w21), .B(w20), .Ci(w16), .S(w10), .Pi(w8), .Gi(w22));   //: @(181, 127) /sz:(64, 63) /sn:0 /p:[ Li0>0 Li1>0 Li2>3 Ro0<1 Ro1<3 Ro2<0 ]
  led g23 (.I(w9));   //: @(233,420) /sn:0 /R:1 /w:[ 0 ] /type:0
  led g24 (.I(w12));   //: @(387,423) /sn:0 /R:2 /w:[ 0 ] /type:0
  CLL g1 (.G0(w34), .P0(w35), .G1(w28), .P1(w29), .G2(w22), .P2(w8), .G3(w3), .P3(w4), .Cin(w14), .C1(w17), .C2(w16), .C3(w0), .C4(w18), .GG(w12), .PG(w9));   //: @(52, 268) /sz:(385, 86) /sn:0 /p:[ Ti0>1 Ti1>7 Ti2>1 Ti3>1 Ti4>1 Ti5>0 Ti6>1 Ti7>1 Ri0>0 To0<0 To1<0 To2<1 Lo0<0 Bo0<1 Bo1<1 ]
  //: dip A (w37) @(-105,62) /w:[ 0 ] /st:3
  //: joint g18 (w16) @(174, 238) /w:[ 1 2 -1 4 ]
  tran g10(.Z(w1), .I(w38[3]));   //: @(-9,70) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  tran g6(.Z(w2), .I(w37[3]));   //: @(29,100) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g7(.Z(w21), .I(w37[2]));   //: @(167,100) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g9(.Z(w33), .I(w37[0]));   //: @(384,100) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  led g22 (.I(w18));   //: @(-23,274) /sn:0 /w:[ 1 ] /type:0
  tran g12(.Z(w26), .I(w38[1]));   //: @(265,70) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  //: dip g5 (w38) @(-44,28) /sn:0 /w:[ 9 ] /st:8
  tran g11(.Z(w20), .I(w38[2]));   //: @(158,70) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  //: switch g14 (w14) @(579,266) /sn:0 /R:1 /w:[ 3 ] /st:0
  //: joint g19 (w8) @(268, 213) /w:[ -1 2 1 4 ]
  led g21 (.I(w11));   //: @(390,-84) /sn:0 /R:3 /w:[ 0 ] /type:2
  concat g20 (.I0(w6), .I1(w7), .I2(w10), .I3(w5), .Z(w11));   //: @(268,-76) /sn:0 /R:1 /w:[ 0 0 0 1 1 ] /dr:0
  PFA g0 (.A(w2), .B(w1), .Ci(w0), .S(w5), .Pi(w4), .Gi(w3));   //: @(62, 126) /sz:(72, 66) /sn:0 /p:[ Li0>0 Li1>0 Li2>0 Ro0<0 Ro1<0 Ro2<0 ]
  //: joint g15 (w14) @(530, 213) /w:[ 2 -1 4 1 ]
  tran g13(.Z(w32), .I(w38[0]));   //: @(376,70) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1

endmodule

module CLA(A, S, B, Cin);
//: interface  /sz:(162, 96) /bd:[ Ti0>A[3:0](24/162) Ti1>B[3:0](61/162) Ri0>Cin(34/96) Bo0<S[3:0](24/162) Bo1<G[3:0](62/162) Bo2<P[3:0](113/162) ]
input [3:0] B;    //: /sn:0 {0}(117,75)(205,75){1}
//: {2}(206,75)(306,75){3}
//: {4}(307,75)(406,75){5}
//: {6}(407,75)(498,75){7}
//: {8}(499,75)(559,75){9}
input [3:0] A;    //: /sn:0 {0}(126,58)(175,58){1}
//: {2}(176,58)(277,58){3}
//: {4}(278,58)(378,58){5}
//: {6}(379,58)(469,58){7}
//: {8}(470,58)(557,58){9}
input Cin;    //: /sn:0 {0}(574,109)(557,109){1}
//: {2}(553,109)(526,109)(526,120){3}
//: {4}(555,111)(555,238)(538,238){5}
output [3:0] S;    //: /sn:0 /dp:1 {0}(639,197)(721,197){1}
wire w16;    //: /sn:0 {0}(412,164)(412,205)(413,205)(413,215){1}
wire w13;    //: /sn:0 {0}(407,122)(407,79){1}
wire w6;    //: /sn:0 {0}(278,123)(278,62){1}
wire w7;    //: /sn:0 {0}(307,123)(307,79){1}
wire w4;    //: /sn:0 {0}(201,164)(201,215){1}
wire w22;    //: /sn:0 {0}(505,165)(505,205)(504,205)(504,215){1}
wire w3;    //: /sn:0 {0}(174,164)(174,182)(633,182){1}
wire w0;    //: /sn:0 {0}(176,122)(176,62){1}
wire w20;    //: /sn:0 /dp:1 {0}(448,215)(448,112)(433,112)(433,122){1}
wire w19;    //: /sn:0 {0}(499,120)(499,79){1}
wire w18;    //: /sn:0 {0}(470,120)(470,62){1}
wire w12;    //: /sn:0 {0}(379,122)(379,62){1}
wire w23;    //: /sn:0 {0}(526,165)(526,205)(527,205)(527,215){1}
wire w10;    //: /sn:0 {0}(313,165)(313,215){1}
wire w21;    //: /sn:0 {0}(478,165)(478,212)(633,212){1}
wire w1;    //: /sn:0 {0}(206,122)(206,79){1}
wire w8;    //: /sn:0 /dp:1 {0}(250,215)(250,112)(234,112)(234,122){1}
wire w17;    //: /sn:0 {0}(433,164)(433,205)(434,205)(434,215){1}
wire w14;    //: /sn:0 /dp:1 {0}(353,215)(353,113)(334,113)(334,123){1}
wire w2;    //: /sn:0 {0}(143,237)(153,237){1}
wire w11;    //: /sn:0 {0}(334,165)(334,205)(335,205)(335,215){1}
wire w15;    //: /sn:0 {0}(386,164)(386,202)(633,202){1}
wire w5;    //: /sn:0 {0}(225,164)(225,205)(226,205)(226,215){1}
wire w9;    //: /sn:0 {0}(286,165)(286,192)(633,192){1}
//: enddecls

  tran g8(.Z(w0), .I(A[3]));   //: @(176,56) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: input g4 (A) @(559,58) /sn:0 /R:2 /w:[ 9 ]
  CLL g16 (.P3(w4), .G3(w5), .P2(w10), .G2(w11), .P1(w16), .G1(w17), .P0(w22), .G0(w23), .Cin(Cin), .C3(w8), .C2(w14), .C1(w20), .C4(w2));   //: @(154, 216) /sz:(383, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>5 To0<0 To1<0 To2<0 Lo0<1 ]
  PFA g3 (.Ci(Cin), .B(w19), .A(w18), .G0(w23), .P0(w22), .S(w21));   //: @(455, 121) /sz:(77, 43) /sn:0 /p:[ Ti0>3 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  concat g17 (.I0(w21), .I1(w15), .I2(w9), .I3(w3), .Z(S));   //: @(638,197) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0
  PFA g2 (.Ci(w20), .B(w13), .A(w12), .G1(w17), .P1(w16), .S(w15));   //: @(364, 123) /sz:(75, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  PFA g1 (.Ci(w14), .B(w7), .A(w6), .G2(w11), .P2(w10), .S(w9));   //: @(263, 124) /sz:(77, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  //: output g18 (S) @(718,197) /sn:0 /w:[ 1 ]
  tran g10(.Z(w19), .I(B[0]));   //: @(499,73) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g6(.Z(w12), .I(A[1]));   //: @(379,56) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g9 (B) @(561,75) /sn:0 /R:2 /w:[ 9 ]
  tran g7(.Z(w6), .I(A[2]));   //: @(278,56) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g12(.Z(w7), .I(B[2]));   //: @(307,73) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: input g14 (Cin) @(576,109) /sn:0 /R:2 /w:[ 0 ]
  tran g11(.Z(w13), .I(B[1]));   //: @(407,73) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g5(.Z(w18), .I(A[0]));   //: @(470,56) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: joint g15 (Cin) @(555, 109) /w:[ 1 -1 2 4 ]
  PFA g0 (.Ci(w8), .B(w1), .A(w0), .G3(w5), .P3(w4), .S(w3));   //: @(160, 123) /sz:(80, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  tran g13(.Z(w1), .I(B[3]));   //: @(206,73) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1

endmodule
