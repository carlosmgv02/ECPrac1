//: version "1.8.7"

module CLL(C1, P3, G3, P0, C3, C4, C0, P1, C2, G0, P2, G2, G1);
//: interface  /sz:(622, 40) /bd:[ Ti0>P3(584/622) Ti1>G3(554/622) Ti2>C3(477/622) Ti3>P2(412/622) Ti4>G2(384/622) Ti5>C2(323/622) Ti6>P1(261/622) Ti7>G1(232/622) Ti8>C1(152/622) Ti9>P0(100/622) Ti10>G0(67/622) Li0>C0(19/40) To0<C0(176/622) Ro0<C4(19/40) ]
input G2;    //: /sn:0 /dp:3 {0}(602,341)(140,341)(140,265)(120,265){1}
//: {2}(116,265)(51,265){3}
//: {4}(118,267)(118,461)(317,461){5}
input C0;    //: /sn:0 {0}(51,65)(205,65){1}
//: {2}(209,65)(401,65)(401,126)(403,126){3}
//: {4}(207,67)(207,155)(241,155){5}
//: {6}(245,155)(278,155)(278,179)(324,179){7}
//: {8}(243,157)(243,250)(249,250){9}
//: {10}(253,250)(326,250){11}
//: {12}(251,252)(251,353)(316,353){13}
input P1;    //: /sn:0 /dp:1 {0}(316,363)(242,363){1}
//: {2}(238,363)(221,363)(221,282){3}
//: {4}(223,280)(326,280){5}
//: {6}(219,280)(210,280)(210,262){7}
//: {8}(212,260)(326,260){9}
//: {10}(208,260)(201,260)(201,211){11}
//: {12}(203,209)(324,209){13}
//: {14}(199,209)(192,209)(192,182){15}
//: {16}(194,180)(264,180)(264,189)(324,189){17}
//: {18}(190,180)(52,180){19}
//: {20}(240,365)(240,399)(316,399){21}
output C3;    //: /sn:0 {0}(661,333)(623,333){1}
input G0;    //: /sn:0 {0}(52,140)(157,140){1}
//: {2}(161,140)(605,140){3}
//: {4}(159,142)(159,204)(168,204){5}
//: {6}(172,204)(324,204){7}
//: {8}(170,206)(170,275)(176,275){9}
//: {10}(180,275)(326,275){11}
//: {12}(178,277)(178,394)(316,394){13}
output C4;    //: /sn:0 /dp:1 {0}(621,423)(658,423){1}
output C2;    //: /sn:0 {0}(660,228)(623,228){1}
input P3;    //: /sn:0 {0}(316,436)(142,436)(142,411){1}
//: {2}(144,409)(316,409){3}
//: {4}(140,409)(109,409)(109,315){5}
//: {6}(111,313)(279,313)(279,373)(316,373){7}
//: {8}(107,313)(49,313){9}
input G1;    //: /sn:0 {0}(602,233)(104,233){1}
//: {2}(100,233)(71,233)(71,202)(51,202){3}
//: {4}(102,235)(102,299)(127,299){5}
//: {6}(131,299)(326,299){7}
//: {8}(129,301)(129,426)(316,426){9}
input G3;    //: /sn:0 /dp:1 {0}(317,466)(100,466)(100,333)(49,333){1}
output C1;    //: /sn:0 {0}(664,138)(626,138){1}
input P0;    //: /sn:0 /dp:1 {0}(52,120)(176,120){1}
//: {2}(180,120)(371,120)(371,131)(403,131){3}
//: {4}(178,122)(178,184)(218,184){5}
//: {6}(222,184)(324,184){7}
//: {8}(220,186)(220,255)(227,255){9}
//: {10}(231,255)(326,255){11}
//: {12}(229,257)(229,358)(316,358){13}
input P2;    //: /sn:0 {0}(316,404)(233,404){1}
//: {2}(229,404)(210,404)(210,370){3}
//: {4}(212,368)(316,368){5}
//: {6}(208,368)(201,368)(201,306){7}
//: {8}(203,304)(326,304){9}
//: {10}(199,304)(185,304)(185,287){11}
//: {12}(187,285)(326,285){13}
//: {14}(183,285)(154,285)(154,245){15}
//: {16}(156,243)(288,243)(288,265)(326,265){17}
//: {18}(152,243)(52,243){19}
//: {20}(231,406)(231,431)(316,431){21}
wire w7;    //: /sn:0 /dp:1 {0}(602,331)(582,331)(582,280)(347,280){1}
wire w4;    //: /sn:0 /dp:1 {0}(602,228)(559,228)(559,207)(345,207){1}
wire w42;    //: /sn:0 {0}(602,336)(574,336)(574,302)(347,302){1}
wire w24;    //: /sn:0 {0}(337,363)(590,363)(590,416)(600,416){1}
wire w8;    //: /sn:0 {0}(424,129)(595,129)(595,135)(605,135){1}
wire w27;    //: /sn:0 {0}(337,401)(584,401)(584,421)(600,421){1}
wire w33;    //: /sn:0 {0}(338,464)(590,464)(590,431)(600,431){1}
wire w2;    //: /sn:0 {0}(345,184)(592,184)(592,223)(602,223){1}
wire w41;    //: /sn:0 {0}(600,426)(572,426)(572,431)(337,431){1}
wire w15;    //: /sn:0 {0}(347,257)(592,257)(592,326)(602,326){1}
//: enddecls

  //: output g4 (C1) @(661,138) /sn:0 /w:[ 0 ]
  and g8 (.I0(C0), .I1(P0), .Z(w8));   //: @(414,129) /sn:0 /w:[ 3 3 0 ]
  //: joint g44 (G0) @(178, 275) /w:[ 10 -1 9 12 ]
  or g3 (.I0(w24), .I1(w27), .I2(w41), .I3(w33), .Z(C4));   //: @(611,423) /sn:0 /w:[ 1 1 0 1 0 ]
  //: input g16 (P3) @(47,313) /sn:0 /w:[ 9 ]
  //: joint g47 (P3) @(109, 313) /w:[ 6 -1 8 5 ]
  //: input g17 (G3) @(47,333) /sn:0 /w:[ 1 ]
  and g26 (.I0(G2), .I1(G3), .Z(w33));   //: @(328,464) /sn:0 /w:[ 5 0 0 ]
  or g2 (.I0(w15), .I1(w7), .I2(w42), .I3(G2), .Z(C3));   //: @(613,333) /sn:0 /w:[ 1 0 0 0 1 ]
  and g23 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .I4(P3), .Z(w24));   //: @(327,363) /sn:0 /w:[ 13 13 0 5 7 0 ]
  //: joint g30 (G0) @(159, 140) /w:[ 2 -1 1 4 ]
  or g1 (.I0(w2), .I1(w4), .I2(G1), .Z(C2));   //: @(613,228) /sn:0 /w:[ 1 0 0 1 ]
  and g24 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w27));   //: @(327,401) /sn:0 /w:[ 13 21 0 3 0 ]
  //: joint g39 (P2) @(185, 285) /w:[ 12 -1 14 11 ]
  //: joint g29 (P0) @(178, 120) /w:[ 2 -1 1 4 ]
  and g18 (.I0(C0), .I1(P0), .I2(P1), .Z(w2));   //: @(335,184) /sn:0 /w:[ 7 7 17 0 ]
  //: input g10 (P0) @(50,120) /sn:0 /w:[ 0 ]
  and g25 (.I0(G1), .I1(P2), .I2(P3), .Z(w41));   //: @(327,431) /sn:0 /w:[ 9 21 0 1 ]
  //: joint g49 (P2) @(231, 404) /w:[ 1 -1 2 20 ]
  //: output g6 (C3) @(658,333) /sn:0 /w:[ 0 ]
  //: joint g50 (P3) @(142, 409) /w:[ 2 -1 4 1 ]
  //: output g7 (C4) @(655,423) /sn:0 /w:[ 1 ]
  //: input g9 (C0) @(49,65) /sn:0 /w:[ 0 ]
  //: joint g35 (G0) @(170, 204) /w:[ 6 -1 5 8 ]
  and g22 (.I0(G1), .I1(P2), .Z(w42));   //: @(337,302) /sn:0 /w:[ 7 9 1 ]
  //: joint g31 (P1) @(192, 180) /w:[ 16 -1 18 15 ]
  //: joint g33 (P0) @(220, 184) /w:[ 6 -1 5 8 ]
  //: joint g36 (P1) @(210, 260) /w:[ 8 -1 10 7 ]
  //: joint g41 (P0) @(229, 255) /w:[ 10 -1 9 12 ]
  //: joint g45 (P1) @(240, 363) /w:[ 1 -1 2 20 ]
  //: joint g40 (C0) @(251, 250) /w:[ 10 -1 9 12 ]
  //: joint g42 (P1) @(221, 280) /w:[ 4 -1 6 3 ]
  //: input g12 (P1) @(50,180) /sn:0 /w:[ 19 ]
  //: joint g28 (C0) @(207, 65) /w:[ 2 -1 1 4 ]
  //: joint g34 (P1) @(201, 209) /w:[ 12 -1 14 11 ]
  //: joint g46 (P2) @(210, 368) /w:[ 4 -1 6 3 ]
  //: output g5 (C2) @(657,228) /sn:0 /w:[ 0 ]
  //: input g11 (G0) @(50,140) /sn:0 /w:[ 0 ]
  //: input g14 (P2) @(50,243) /sn:0 /w:[ 19 ]
  and g19 (.I0(G0), .I1(P1), .Z(w4));   //: @(335,207) /sn:0 /w:[ 7 13 1 ]
  and g21 (.I0(G0), .I1(P1), .I2(P2), .Z(w7));   //: @(337,280) /sn:0 /w:[ 11 5 13 1 ]
  and g20 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .Z(w15));   //: @(337,257) /sn:0 /w:[ 11 11 9 17 0 ]
  //: joint g32 (C0) @(243, 155) /w:[ 6 -1 5 8 ]
  or g0 (.I0(w8), .I1(G0), .Z(C1));   //: @(616,138) /sn:0 /w:[ 1 3 1 ]
  //: input g15 (G2) @(49,265) /sn:0 /w:[ 3 ]
  //: joint g38 (G1) @(102, 233) /w:[ 1 -1 2 4 ]
  //: joint g43 (P2) @(201, 304) /w:[ 8 -1 10 7 ]
  //: joint g27 (G2) @(118, 265) /w:[ 1 -1 2 4 ]
  //: joint g48 (G1) @(129, 299) /w:[ 6 -1 5 8 ]
  //: joint g37 (P2) @(154, 243) /w:[ 16 -1 18 15 ]
  //: input g13 (G1) @(49,202) /sn:0 /w:[ 3 ]

endmodule

module PFA(Pi, A, Ci, Gi, S, B);
//: interface  /sz:(100, 97) /bd:[ Ti0>A(14/100) Ti1>B(50/100) Li0>Ci(46/97) Bo0<Gi(61/100) Ro0<S(32/97) Ro1<Pi(67/97) ]
input B;    //: /sn:0 {0}(184,223)(195,223){1}
//: {2}(199,223)(226,223)(226,207)(234,207){3}
//: {4}(197,225)(197,256){5}
//: {6}(199,258)(308,258){7}
//: {8}(197,260)(197,293)(309,293){9}
output Gi;    //: /sn:0 /dp:1 {0}(330,291)(354,291){1}
input A;    //: /sn:0 {0}(186,202)(214,202){1}
//: {2}(218,202)(234,202){3}
//: {4}(216,204)(216,251){5}
//: {6}(218,253)(308,253){7}
//: {8}(216,255)(216,288)(309,288){9}
output Pi;    //: /sn:0 /dp:1 {0}(329,256)(351,256){1}
input Ci;    //: /sn:0 /dp:1 {0}(305,227)(274,227)(274,241)(187,241){1}
output S;    //: /sn:0 {0}(358,225)(326,225){1}
wire w11;    //: /sn:0 {0}(255,205)(295,205)(295,222)(305,222){1}
//: enddecls

  //: output g8 (Pi) @(348,256) /sn:0 /w:[ 1 ]
  //: input g4 (A) @(184,202) /sn:0 /w:[ 0 ]
  xor g3 (.I0(A), .I1(B), .Z(w11));   //: @(245,205) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  xor g2 (.I0(w11), .I1(Ci), .Z(S));   //: @(316,225) /sn:0 /delay:" 2" /w:[ 1 0 1 ]
  or g1 (.I0(A), .I1(B), .Z(Pi));   //: @(319,256) /sn:0 /w:[ 7 7 0 ]
  //: joint g10 (A) @(216, 202) /w:[ 2 -1 1 4 ]
  //: input g6 (Ci) @(185,241) /sn:0 /w:[ 1 ]
  //: output g9 (Gi) @(351,291) /sn:0 /w:[ 1 ]
  //: output g7 (S) @(355,225) /sn:0 /w:[ 0 ]
  //: joint g12 (A) @(216, 253) /w:[ 6 5 -1 8 ]
  //: joint g11 (B) @(197, 223) /w:[ 2 -1 1 4 ]
  //: input g5 (B) @(182,223) /sn:0 /w:[ 0 ]
  and g0 (.I0(A), .I1(B), .Z(Gi));   //: @(320,291) /sn:0 /w:[ 9 9 0 ]
  //: joint g13 (B) @(197, 258) /w:[ 6 5 -1 8 ]

endmodule

module CLA16(A, Cout, S, B, Cin);
//: interface  /sz:(214, 188) /bd:[ Ti0>B[15:0](126/214) Ti1>A[15:0](46/214) Li0>Cin(64/188) Bo0<S[15:0](134/214) Ro0<Cout(74/188) ]
input [15:0] B;    //: /sn:0 {0}(-300,-257)(-177,-257){1}
//: {2}(-176,-257)(-30,-257){3}
//: {4}(-29,-257)(138,-257){5}
//: {6}(139,-257)(307,-257){7}
//: {8}(308,-257)(427,-257){9}
input [15:0] A;    //: /sn:0 {0}(-298,-282)(-242,-282){1}
//: {2}(-241,-282)(-95,-282){3}
//: {4}(-94,-282)(73,-282){5}
//: {6}(74,-282)(242,-282){7}
//: {8}(243,-282)(427,-282){9}
input Cin;    //: /sn:0 {0}(-295,-154)(-265,-154){1}
output Cout;    //: /sn:0 {0}(385,245)(343,245){1}
output [15:0] S;    //: /sn:0 {0}(512,356)(553,356){1}
wire [3:0] w13;    //: /sn:0 {0}(117,155)(117,351)(506,351){1}
wire [3:0] w16;    //: /sn:0 {0}(243,192)(243,-278){1}
wire [3:0] w6;    //: /sn:0 {0}(-94,-63)(-94,-278){1}
wire w4;    //: /sn:0 {0}(-141,-148)(-128,-148)(-128,-16)(-118,-16){1}
wire [3:0] w0;    //: /sn:0 {0}(-176,-201)(-176,-253){1}
wire [3:0] w3;    //: /sn:0 {0}(-198,-101)(-198,371)(506,371){1}
wire [3:0] w18;    //: /sn:0 {0}(286,292)(286,341)(506,341){1}
wire [3:0] w10;    //: /sn:0 {0}(139,55)(139,-253){1}
wire [3:0] w1;    //: /sn:0 {0}(-241,-201)(-241,-278){1}
wire [3:0] w8;    //: /sn:0 {0}(-51,37)(-51,361)(506,361){1}
wire w14;    //: /sn:0 {0}(174,108)(209,108)(209,239)(219,239){1}
wire [3:0] w11;    //: /sn:0 {0}(74,55)(74,-278){1}
wire [3:0] w15;    //: /sn:0 {0}(308,192)(308,-253){1}
wire [3:0] w5;    //: /sn:0 {0}(-29,-63)(-29,-253){1}
wire w9;    //: /sn:0 {0}(6,-10)(40,-10)(40,102)(50,102){1}
//: enddecls

  tran g8(.Z(w6), .I(A[7:4]));   //: @(-94,-284) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: input g4 (A) @(-300,-282) /sn:0 /w:[ 0 ]
  //: output g16 (Cout) @(382,245) /sn:0 /w:[ 0 ]
  CLA g3 (.A(w16), .B(w15), .C0(w14), .S(w18), .C4(Cout));   //: @(220, 193) /sz:(122, 98) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<1 ]
  concat g17 (.I0(w3), .I1(w8), .I2(w13), .I3(w18), .Z(S));   //: @(511,356) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0
  CLA g2 (.A(w11), .B(w10), .C0(w9), .S(w13), .C4(w14));   //: @(51, 56) /sz:(122, 98) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<0 ]
  CLA g1 (.A(w6), .B(w5), .C0(w4), .S(w8), .C4(w9));   //: @(-117, -62) /sz:(122, 98) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<0 ]
  tran g10(.Z(w11), .I(A[11:8]));   //: @(74,-284) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g6(.Z(w1), .I(A[3:0]));   //: @(-241,-284) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g9(.Z(w5), .I(B[7:4]));   //: @(-29,-259) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g7(.Z(w0), .I(B[3:0]));   //: @(-176,-259) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g12(.Z(w16), .I(A[15:12]));   //: @(243,-284) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: output g14 (S) @(550,356) /sn:0 /w:[ 1 ]
  tran g11(.Z(w10), .I(B[11:8]));   //: @(139,-259) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g5 (B) @(-302,-257) /sn:0 /w:[ 0 ]
  //: input g15 (Cin) @(-297,-154) /sn:0 /w:[ 0 ]
  CLA g0 (.A(w1), .B(w0), .C0(Cin), .S(w3), .C4(w4));   //: @(-264, -200) /sz:(122, 98) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<0 ]
  tran g13(.Z(w15), .I(B[15:12]));   //: @(308,-259) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1

endmodule

module main;    //: root_module
wire w13;    //: /sn:0 {0}(43,174)(9,174)(9,287)(-65,287){1}
wire w65;    //: /sn:0 {0}(43,124)(-55,124)(-55,143)(-65,143){1}
wire w7;    //: /sn:0 /dp:1 {0}(43,184)(-49,184)(-49,316)(-65,316){1}
wire w88;    //: /sn:0 {0}(426,280)(382,280)(382,183)(320,183){1}
wire w81;    //: /sn:0 {0}(-64,113)(18,113)(18,114)(43,114){1}
wire w72;    //: /sn:0 {0}(320,113)(402,113)(402,75)(427,75){1}
wire w62;    //: /sn:0 {0}(43,154)(-8,154)(-8,230)(-65,230){1}
wire w82;    //: /sn:0 {0}(426,309)(376,309)(376,193)(320,193){1}
wire w3;    //: /sn:0 /dp:1 {0}(43,194)(-58,194)(-58,345)(-65,345){1}
wire [3:0] w60;    //: /sn:0 {0}(438,406)(438,471)(313,471){1}
wire w71;    //: /sn:0 {0}(320,103)(384,103)(384,46)(427,46){1}
wire w73;    //: /sn:0 {0}(320,123)(417,123)(417,104)(427,104){1}
wire w66;    //: /sn:0 {0}(320,53)(420,53)(420,-98)(427,-98){1}
wire w18;    //: /sn:0 {0}(43,164)(0,164)(0,258)(-65,258){1}
wire [15:0] w10;    //: /sn:0 /dp:1 {0}(49,119)(109,119)(109,162)(135,162)(135,213){1}
wire w63;    //: /sn:0 {0}(43,144)(-22,144)(-22,201)(-65,201){1}
wire w70;    //: /sn:0 {0}(320,73)(353,73)(353,-40)(427,-40){1}
wire w84;    //: /sn:0 {0}(426,221)(402,221)(402,163)(320,163){1}
wire w86;    //: /sn:0 {0}(426,192)(407,192)(407,153)(320,153){1}
wire w68;    //: /sn:0 {0}(320,83)(362,83)(362,-11)(427,-11){1}
wire [3:0] w32;    //: /sn:0 {0}(353,405)(353,441)(313,441){1}
wire w8;    //: /sn:0 {0}(66,278)(88,278){1}
wire w89;    //: /sn:0 {0}(426,338)(367,338)(367,203)(320,203){1}
wire w75;    //: /sn:0 {0}(-64,-62)(-14,-62)(-14,54)(43,54){1}
wire w67;    //: /sn:0 {0}(320,93)(370,93)(370,17)(427,17){1}
wire w80;    //: /sn:0 {0}(-64,84)(-56,84)(-56,104)(43,104){1}
wire [3:0] w33;    //: /sn:0 {0}(384,405)(384,451)(313,451){1}
wire w69;    //: /sn:0 {0}(320,63)(411,63)(411,-69)(427,-69){1}
wire w78;    //: /sn:0 {0}(-64,55)(-45,55)(-45,94)(43,94){1}
wire w74;    //: /sn:0 {0}(-64,-91)(-5,-91)(-5,44)(43,44){1}
wire [15:0] w90;    //: /sn:0 {0}(314,128)(215,128)(215,213){1}
wire w85;    //: /sn:0 {0}(426,134)(344,134)(344,133)(320,133){1}
wire w83;    //: /sn:0 {0}(426,163)(418,163)(418,143)(320,143){1}
wire [3:0] w61;    //: /sn:0 {0}(411,406)(411,461)(313,461){1}
wire w87;    //: /sn:0 {0}(426,251)(393,251)(393,173)(320,173){1}
wire w64;    //: /sn:0 {0}(43,134)(-40,134)(-40,172)(-65,172){1}
wire [15:0] S;    //: /sn:0 {0}(307,456)(223,456)(223,403){1}
wire w76;    //: /sn:0 {0}(-64,-33)(-20,-33)(-20,64)(43,64){1}
wire w9;    //: /sn:0 /dp:1 {0}(329,288)(304,288){1}
wire w79;    //: /sn:0 {0}(-64,26)(-40,26)(-40,84)(43,84){1}
wire w77;    //: /sn:0 {0}(-64,-4)(-31,-4)(-31,74)(43,74){1}
//: enddecls

  //: switch g75 (w66) @(445,-98) /sn:0 /R:2 /w:[ 1 ] /st:1
  led g4 (.I(w32));   //: @(353,398) /sn:0 /w:[ 0 ] /type:1
  concat g3 (.I0(w32), .I1(w33), .I2(w61), .I3(w60), .Z(S));   //: @(308,456) /sn:0 /R:2 /w:[ 1 1 1 1 0 ] /dr:0
  //: switch g90 (w86) @(444,192) /sn:0 /R:2 /w:[ 0 ] /st:1
  //: switch g2 (w8) @(49,278) /sn:0 /w:[ 0 ] /st:1
  //: switch g91 (w87) @(444,251) /sn:0 /R:2 /w:[ 0 ] /st:1
  //: switch g74 (w3) @(-82,345) /sn:0 /w:[ 1 ] /st:1
  //: switch g86 (w72) @(445,75) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: switch g77 (w67) @(445,17) /sn:0 /R:2 /w:[ 1 ] /st:1
  led g1 (.I(w9));   //: @(336,288) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: switch g60 (w75) @(-81,-62) /sn:0 /w:[ 0 ] /st:1
  //: switch g82 (w73) @(445,104) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: switch g70 (w62) @(-82,230) /sn:0 /w:[ 1 ] /st:1
  //: switch g65 (w80) @(-81,84) /sn:0 /w:[ 0 ] /st:1
  //: switch g64 (w79) @(-81,26) /sn:0 /w:[ 0 ] /st:1
  //: switch g72 (w18) @(-82,258) /sn:0 /w:[ 1 ] /st:1
  //: switch g73 (w7) @(-82,316) /sn:0 /w:[ 1 ] /st:1
  //: switch g68 (w65) @(-82,143) /sn:0 /w:[ 1 ] /st:1
  concat g58 (.I0(w3), .I1(w7), .I2(w13), .I3(w18), .I4(w62), .I5(w63), .I6(w64), .I7(w65), .I8(w81), .I9(w80), .I10(w78), .I11(w79), .I12(w77), .I13(w76), .I14(w75), .I15(w74), .Z(w10));   //: @(48,119) /sn:0 /w:[ 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 ] /dr:0
  led g56 (.I(w60));   //: @(438,399) /sn:0 /w:[ 0 ] /type:1
  //: switch g71 (w13) @(-82,287) /sn:0 /w:[ 1 ] /st:1
  //: switch g59 (w74) @(-81,-91) /sn:0 /w:[ 0 ] /st:1
  //: switch g87 (w71) @(445,46) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: switch g85 (w70) @(445,-40) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: switch g67 (w64) @(-82,172) /sn:0 /w:[ 1 ] /st:1
  //: switch g83 (w69) @(445,-69) /sn:0 /R:2 /w:[ 1 ] /st:1
  concat g81 (.I0(w66), .I1(w69), .I2(w70), .I3(w68), .I4(w67), .I5(w71), .I6(w72), .I7(w73), .I8(w85), .I9(w83), .I10(w86), .I11(w84), .I12(w87), .I13(w88), .I14(w82), .I15(w89), .Z(w90));   //: @(315,128) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 ] /dr:0
  //: switch g69 (w63) @(-82,201) /sn:0 /w:[ 1 ] /st:1
  //: switch g66 (w81) @(-81,113) /sn:0 /w:[ 0 ] /st:1
  led g57 (.I(w61));   //: @(411,399) /sn:0 /w:[ 0 ] /type:1
  //: switch g84 (w89) @(444,338) /sn:0 /R:2 /w:[ 0 ] /st:1
  led g5 (.I(w33));   //: @(384,398) /sn:0 /w:[ 0 ] /type:1
  //: switch g61 (w76) @(-81,-33) /sn:0 /w:[ 0 ] /st:1
  //: switch g79 (w84) @(444,221) /sn:0 /R:2 /w:[ 0 ] /st:1
  //: switch g78 (w83) @(444,163) /sn:0 /R:2 /w:[ 0 ] /st:1
  //: switch g63 (w78) @(-81,55) /sn:0 /w:[ 0 ] /st:1
  //: switch g89 (w88) @(444,280) /sn:0 /R:2 /w:[ 0 ] /st:1
  CLA16 g0 (.A(w10), .B(w90), .Cin(w8), .S(S), .Cout(w9));   //: @(89, 214) /sz:(214, 188) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Ro0<1 ]
  //: switch g62 (w77) @(-81,-4) /sn:0 /w:[ 0 ] /st:1
  //: switch g88 (w85) @(444,134) /sn:0 /R:2 /w:[ 0 ] /st:1
  //: switch g80 (w68) @(445,-11) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: switch g76 (w82) @(444,309) /sn:0 /R:2 /w:[ 0 ] /st:1

endmodule

module CLA(A, C4, B, S, C0);
//: interface  /sz:(122, 98) /bd:[ Ti0>B[3:0](88/122) Ti1>A[3:0](23/122) Li0>C0(46/98) Bo0<S[3:0](66/122) Ro0<C4(52/98) ]
input [3:0] B;    //: /sn:0 /dp:1 {0}(40,86)(137,86){1}
//: {2}(138,86)(301,86){3}
//: {4}(302,86)(459,86){5}
//: {6}(460,86)(621,86){7}
//: {8}(622,86)(726,86){9}
input C0;    //: /sn:0 {0}(30,251)(40,251){1}
//: {2}(44,251)(52,251)(52,215)(87,215){3}
//: {4}(42,253)(42,372)(61,372){5}
input [3:0] A;    //: /sn:0 {0}(42,61)(101,61){1}
//: {2}(102,61)(138,61)(138,61)(265,61){3}
//: {4}(266,61)(423,61){5}
//: {6}(424,61)(585,61){7}
//: {8}(586,61)(732,61){9}
output C4;    //: /sn:0 {0}(739,372)(685,372){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(760,529)(739,529){1}
wire w6;    //: /sn:0 {0}(302,170)(302,90){1}
wire w13;    //: /sn:0 {0}(424,170)(424,65){1}
wire w7;    //: /sn:0 {0}(266,170)(266,65){1}
wire w34;    //: /sn:0 /dp:1 {0}(549,352)(549,220)(571,220){1}
wire w0;    //: /sn:0 {0}(138,168)(138,90){1}
wire w3;    //: /sn:0 /dp:1 {0}(733,534)(381,534)(381,203)(353,203){1}
wire w29;    //: /sn:0 /dp:1 {0}(321,352)(321,294)(368,294)(368,238)(353,238){1}
wire w12;    //: /sn:0 {0}(460,170)(460,90){1}
wire w18;    //: /sn:0 {0}(622,173)(622,90){1}
wire w19;    //: /sn:0 {0}(586,173)(586,65){1}
wire w10;    //: /sn:0 {0}(733,514)(705,514)(705,206)(673,206){1}
wire w21;    //: /sn:0 {0}(595,272)(595,352){1}
wire w1;    //: /sn:0 {0}(102,168)(102,65){1}
wire w31;    //: /sn:0 /dp:1 {0}(385,352)(385,217)(409,217){1}
wire w32;    //: /sn:0 /dp:1 {0}(471,352)(471,296)(525,296)(525,244)(511,244){1}
wire w8;    //: /sn:0 {0}(733,524)(541,524)(541,218)(511,218){1}
wire w27;    //: /sn:0 /dp:1 {0}(112,352)(112,267){1}
wire w35;    //: /sn:0 /dp:1 {0}(638,352)(638,301)(688,301)(688,241)(673,241){1}
wire w28;    //: /sn:0 {0}(229,352)(229,217)(251,217){1}
wire w2;    //: /sn:0 {0}(733,544)(212,544)(212,201)(189,201){1}
wire w15;    //: /sn:0 {0}(433,269)(433,352){1}
wire w9;    //: /sn:0 {0}(278,269)(278,352){1}
wire w26;    //: /sn:0 /dp:1 {0}(137,352)(137,320)(201,320)(201,236)(189,236){1}
//: enddecls

  //: input g4 (A) @(40,61) /sn:0 /w:[ 0 ]
  tran g8(.Z(w7), .I(A[1]));   //: @(266,59) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  PFA g3 (.A(w19), .B(w18), .Ci(w34), .Gi(w21), .S(w10), .Pi(w35));   //: @(572, 174) /sz:(100, 97) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<1 Ro1<1 ]
  //: joint g16 (C0) @(42, 251) /w:[ 2 -1 1 4 ]
  //: output g17 (C4) @(736,372) /sn:0 /w:[ 0 ]
  PFA g2 (.A(w13), .B(w12), .Ci(w31), .Gi(w15), .S(w8), .Pi(w32));   //: @(410, 171) /sz:(100, 97) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<1 Ro1<1 ]
  PFA g1 (.A(w7), .B(w6), .Ci(w28), .Gi(w9), .S(w3), .Pi(w29));   //: @(252, 171) /sz:(100, 97) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<1 Ro1<1 ]
  concat g18 (.I0(w2), .I1(w3), .I2(w8), .I3(w10), .Z(S));   //: @(738,529) /sn:0 /w:[ 0 0 0 0 1 ] /dr:0
  tran g10(.Z(w13), .I(A[2]));   //: @(424,59) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g6(.Z(w1), .I(A[0]));   //: @(102,59) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g9(.Z(w6), .I(B[1]));   //: @(302,84) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g7(.Z(w0), .I(B[0]));   //: @(138,84) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g12(.Z(w19), .I(A[3]));   //: @(586,59) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: input g5 (B) @(38,86) /sn:0 /w:[ 0 ]
  tran g11(.Z(w12), .I(B[2]));   //: @(460,84) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  CLL g14 (.P3(w21), .G3(w35), .P2(w15), .G2(w32), .P1(w9), .G1(w29), .P0(w27), .G0(w26), .C0(C0), .C3(w34), .C2(w31), .C1(w28), .C4(C4));   //: @(62, 353) /sz:(622, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>1 Ti3>0 Ti4>1 Ti5>0 Ti6>0 Ti7>0 Li0>5 To0<0 To1<0 To2<0 Ro0<1 ]
  //: output g19 (S) @(757,529) /sn:0 /w:[ 0 ]
  PFA g0 (.A(w1), .B(w0), .Ci(C0), .Gi(w27), .S(w2), .Pi(w26));   //: @(88, 169) /sz:(100, 97) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>3 Bo0<1 Ro0<1 Ro1<1 ]
  //: input g15 (C0) @(28,251) /sn:0 /w:[ 0 ]
  tran g13(.Z(w18), .I(B[3]));   //: @(622,84) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1

endmodule
