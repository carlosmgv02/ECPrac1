//: version "1.8.7"

module FA(Cout, S, Cin, B, A);
//: interface  /sz:(225, 114) /bd:[ Ti0>B(166/225) Ti1>A(36/225) Ri0>Cin(52/114) Lo0<Cout(58/114) Bo0<S(117/225) ]
input B;    //: /sn:0 {0}(143,173)(159,173){1}
//: {2}(163,173)(176,173)(176,104)(186,104){3}
//: {4}(161,175)(161,176)(242,176)(242,152)(252,152){5}
input A;    //: /sn:0 {0}(130,98)(150,98){1}
//: {2}(154,98)(176,98)(176,99)(186,99){3}
//: {4}(152,100)(152,147)(252,147){5}
input Cin;    //: /sn:0 {0}(143,199)(213,199)(213,125){1}
//: {2}(215,123)(225,123)(225,124)(253,124){3}
//: {4}(213,121)(213,107)(223,107){5}
output Cout;    //: /sn:0 /dp:1 {0}(324,137)(347,137)(347,136)(357,136){1}
output S;    //: /sn:0 /dp:1 {0}(244,105)(348,105){1}
wire w4;    //: /sn:0 {0}(274,127)(293,127)(293,134)(303,134){1}
wire w2;    //: /sn:0 {0}(207,102)(215,102){1}
//: {2}(219,102)(223,102){3}
//: {4}(217,104)(217,129)(253,129){5}
wire w5;    //: /sn:0 {0}(273,150)(293,150)(293,139)(303,139){1}
//: enddecls

  //: joint g8 (Cin) @(213, 123) /w:[ 2 4 -1 1 ]
  //: output g4 (Cout) @(354,136) /sn:0 /w:[ 1 ]
  //: output g3 (S) @(345,105) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(141,199) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(141,173) /sn:0 /w:[ 0 ]
  and g10 (.I0(A), .I1(B), .Z(w5));   //: @(263,150) /sn:0 /tech:unit /w:[ 5 5 0 ]
  xor g6 (.I0(w2), .I1(Cin), .Z(S));   //: @(234,105) /sn:0 /delay:" 2" /w:[ 3 5 0 ]
  //: joint g9 (w2) @(217, 102) /w:[ 2 -1 1 4 ]
  and g7 (.I0(Cin), .I1(w2), .Z(w4));   //: @(264,127) /sn:0 /tech:unit /w:[ 3 5 0 ]
  //: joint g12 (B) @(161, 173) /w:[ 2 -1 1 4 ]
  //: joint g11 (A) @(152, 98) /w:[ 2 -1 1 4 ]
  xor g5 (.I0(A), .I1(B), .Z(w2));   //: @(197,102) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  //: input g0 (A) @(128,98) /sn:0 /w:[ 0 ]
  or g13 (.I0(w4), .I1(w5), .Z(Cout));   //: @(314,137) /sn:0 /tech:unit /w:[ 1 1 0 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(95,193)(164,193)(164,159)(174,159){1}
wire w7;    //: /sn:0 {0}(111,275)(164,275)(164,196)(174,196){1}
wire w4;    //: /sn:0 {0}(322,174)(344,174)(344,199)(359,199)(359,189){1}
wire w3;    //: /sn:0 {0}(322,123)(384,123)(384,114){1}
wire w5;    //: /sn:0 {0}(108,128)(164,128)(164,124)(174,124){1}
//: enddecls

  led g4 (.I(w3));   //: @(384,107) /sn:0 /w:[ 1 ] /type:0
  //: switch g3 (w7) @(94,275) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w6) @(78,193) /sn:0 /w:[ 0 ] /st:0
  //: switch g1 (w5) @(91,128) /sn:0 /w:[ 0 ] /st:0
  led g5 (.I(w4));   //: @(359,182) /sn:0 /w:[ 1 ] /type:0
  FA g0 (.Cin(w7), .B(w6), .A(w5), .Cout(w4), .S(w3));   //: @(175, 101) /sz:(146, 136) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Ro0<0 Ro1<0 ]

endmodule
