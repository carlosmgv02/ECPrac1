//: version "1.8.7"

module FullAdder2(A, Cin, B, Cout, S);
//: interface  /sz:(96, 63) /bd:[ Ti0>B(51/96) Ti1>A(14/96) Li0>Cin(26/63) Bo0<S(61/96) Bo1<Cout(28/96) ]
input B;    //: /sn:0 /dp:1 {0}(198,211)(186,211){1}
//: {2}(182,211)(159,211)(159,239){3}
//: {4}(157,241)(139,241){5}
//: {6}(159,243)(159,330)(199,330){7}
//: {8}(184,213)(184,305)(198,305){9}
input A;    //: /sn:0 {0}(136,206)(150,206){1}
//: {2}(154,206)(165,206){3}
//: {4}(169,206)(198,206){5}
//: {6}(167,208)(167,271)(198,271){7}
//: {8}(152,208)(152,300)(198,300){9}
input Cin;    //: /sn:0 {0}(143,304)(171,304){1}
//: {2}(173,302)(173,278){3}
//: {4}(175,276)(198,276){5}
//: {6}(173,274)(173,225)(281,225){7}
//: {8}(173,306)(173,335)(199,335){9}
output Cout;    //: /sn:0 {0}(412,321)(386,321){1}
output S;    //: /sn:0 /dp:1 {0}(302,223)(352,223){1}
wire w8;    //: /sn:0 {0}(219,274)(275,274)(275,287)(285,287){1}
wire w17;    //: /sn:0 {0}(306,290)(355,290)(355,318)(365,318){1}
wire w14;    //: /sn:0 {0}(220,333)(355,333)(355,323)(365,323){1}
wire w2;    //: /sn:0 {0}(219,209)(271,209)(271,220)(281,220){1}
wire w11;    //: /sn:0 {0}(219,303)(275,303)(275,292)(285,292){1}
//: enddecls

  and g4 (.I0(B), .I1(Cin), .Z(w14));   //: @(210,333) /sn:0 /w:[ 7 9 0 ]
  //: input g8 (A) @(134,206) /sn:0 /w:[ 0 ]
  and g3 (.I0(A), .I1(B), .Z(w11));   //: @(209,303) /sn:0 /w:[ 9 9 0 ]
  //: joint g16 (A) @(152, 206) /w:[ 2 -1 1 8 ]
  //: joint g17 (B) @(184, 211) /w:[ 1 -1 2 8 ]
  and g2 (.I0(A), .I1(Cin), .Z(w8));   //: @(209,274) /sn:0 /w:[ 7 5 0 ]
  xor g1 (.I0(w2), .I1(Cin), .Z(S));   //: @(292,223) /sn:0 /delay:" 2" /w:[ 1 7 0 ]
  //: input g10 (Cin) @(141,304) /sn:0 /w:[ 0 ]
  or g6 (.I0(w17), .I1(w14), .Z(Cout));   //: @(376,321) /sn:0 /w:[ 1 1 1 ]
  //: joint g7 (A) @(167, 206) /w:[ 4 -1 3 6 ]
  //: input g9 (B) @(137,241) /sn:0 /w:[ 5 ]
  //: output g12 (Cout) @(409,321) /sn:0 /w:[ 0 ]
  or g5 (.I0(w8), .I1(w11), .Z(w17));   //: @(296,290) /sn:0 /w:[ 1 1 0 ]
  //: output g11 (S) @(349,223) /sn:0 /w:[ 1 ]
  //: joint g14 (Cin) @(173, 276) /w:[ 4 6 -1 3 ]
  xor g0 (.I0(A), .I1(B), .Z(w2));   //: @(209,209) /sn:0 /delay:" 2" /w:[ 5 0 0 ]
  //: joint g15 (Cin) @(173, 304) /w:[ -1 2 1 8 ]
  //: joint g13 (B) @(159, 241) /w:[ -1 3 4 6 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(341,136)(344,136)(344,203){1}
wire w0;    //: /sn:0 {0}(257,230)(292,230){1}
wire w1;    //: /sn:0 {0}(321,287)(321,268){1}
wire w2;    //: /sn:0 {0}(354,287)(354,268){1}
wire w5;    //: /sn:0 {0}(294,169)(307,169)(307,203){1}
//: enddecls

  led g4 (.I(w1));   //: @(321,294) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: switch g3 (w0) @(240,230) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w6) @(324,136) /sn:0 /w:[ 0 ] /st:0
  //: switch g1 (w5) @(277,169) /sn:0 /w:[ 0 ] /st:0
  led g5 (.I(w2));   //: @(354,294) /sn:0 /R:2 /w:[ 0 ] /type:0
  FullAdder2 g0 (.B(w6), .A(w5), .Cin(w0), .S(w2), .Cout(w1));   //: @(293, 204) /sz:(96, 63) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Bo1<1 ]

endmodule
