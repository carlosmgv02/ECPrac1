//: version "1.8.7"

module CPA16(Cout, Cin, B, A, S);
//: interface  /sz:(144, 70) /bd:[ Ti0>B[15:0](98/144) Ti1>A[15:0](32/144) Li0>Cin(41/70) Bo0<S[15:0](95/144) Bo1<Cout(46/144) ]
input [15:0] B;    //: /sn:0 {0}(39,-32)(98,-32){1}
//: {2}(99,-32)(111,-32){3}
//: {4}(112,-32)(129,-32){5}
//: {6}(130,-32)(146,-32){7}
//: {8}(147,-32)(274,-32){9}
//: {10}(275,-32)(293,-32){11}
//: {12}(294,-32)(313,-32){13}
//: {14}(314,-32)(330,-32){15}
//: {16}(331,-32)(520,-32){17}
//: {18}(521,-32)(535,-32){19}
//: {20}(536,-32)(552,-32){21}
//: {22}(553,-32)(569,-32){23}
//: {24}(570,-32)(729,-32){25}
//: {26}(730,-32)(746,-32){27}
//: {28}(747,-32)(762,-32){29}
//: {30}(763,-32)(782,-32){31}
//: {32}(783,-32)(832,-32){33}
input [15:0] A;    //: /sn:0 {0}(39,73)(83,73){1}
//: {2}(84,73)(100,73){3}
//: {4}(101,73)(124,73){5}
//: {6}(125,73)(143,73){7}
//: {8}(144,73)(367,73){9}
//: {10}(368,73)(388,73){11}
//: {12}(389,73)(407,73){13}
//: {14}(408,73)(424,73){15}
//: {16}(425,73)(540,73){17}
//: {18}(541,73)(557,73){19}
//: {20}(558,73)(579,73){21}
//: {22}(580,73)(596,73){23}
//: {24}(597,73)(724,73){25}
//: {26}(725,73)(742,73){27}
//: {28}(743,73)(760,73){29}
//: {30}(761,73)(777,73){31}
//: {32}(778,73)(820,73){33}
input Cin;    //: /sn:0 {0}(321,234)(321,281)(180,281){1}
output Cout;    //: /sn:0 /dp:1 {0}(803,236)(803,261)(931,261){1}
output [15:0] S;    //: /sn:0 /dp:1 {0}(958,359)(1002,359){1}
wire w16;    //: /sn:0 {0}(497,234)(497,259)(272,259)(272,234){1}
wire w13;    //: /sn:0 {0}(449,96)(425,96)(425,77){1}
wire w6;    //: /sn:0 {0}(101,77)(101,123)(161,123){1}
wire w58;    //: /sn:0 {0}(952,334)(714,334)(714,319){1}
wire w7;    //: /sn:0 {0}(368,77)(368,126)(449,126){1}
wire w50;    //: /sn:0 {0}(952,414)(353,414)(353,377){1}
wire w34;    //: /sn:0 {0}(588,-2)(553,-2)(553,-28){1}
wire w59;    //: /sn:0 {0}(952,324)(737,324)(737,319){1}
wire w62;    //: /sn:0 {0}(952,294)(887,294)(887,280){1}
wire w39;    //: /sn:0 {0}(612,95)(597,95)(597,77){1}
wire [3:0] w25;    //: /sn:0 /dp:1 {0}(361,2)(499,2)(499,188){1}
wire [3:0] w4;    //: /sn:0 {0}(300,234)(300,373)(313,373){1}
//: {2}(314,373)(322,373)(322,373)(333,373){3}
//: {4}(334,373)(352,373){5}
//: {6}(353,373)(370,373){7}
//: {8}(371,373)(381,373){9}
wire w56;    //: /sn:0 {0}(952,354)(676,354)(676,319){1}
wire w3;    //: /sn:0 {0}(747,-28)(747,7)(796,7){1}
wire w36;    //: /sn:0 {0}(558,77)(558,115)(612,115){1}
wire w0;    //: /sn:0 {0}(541,77)(541,125)(612,125){1}
wire w22;    //: /sn:0 {0}(168,-14)(147,-14)(147,-28){1}
wire w60;    //: /sn:0 {0}(952,314)(839,314)(839,280){1}
wire [3:0] w20;    //: /sn:0 /dp:1 {0}(174,1)(323,1)(323,188){1}
wire w29;    //: /sn:0 {0}(796,-3)(763,-3)(763,-28){1}
wire [3:0] w30;    //: /sn:0 {0}(666,238)(666,315)(675,315){1}
//: {2}(676,315)(691,315){3}
//: {4}(692,315)(713,315){5}
//: {6}(714,315)(736,315){7}
//: {8}(737,315)(759,315){9}
wire w42;    //: /sn:0 {0}(334,377)(334,424)(952,424){1}
wire [3:0] w37;    //: /sn:0 /dp:1 {0}(618,110)(641,110)(641,192){1}
wire w19;    //: /sn:0 {0}(112,-28)(112,6)(168,6){1}
wire [3:0] w18;    //: /sn:0 {0}(557,338)(545,338){1}
//: {2}(544,338)(530,338)(530,339)(517,339){3}
//: {4}(516,339)(495,339){5}
//: {6}(494,339)(481,339){7}
//: {8}(480,339)(476,339)(476,234){9}
wire w12;    //: /sn:0 {0}(449,106)(408,106)(408,77){1}
wire w63;    //: /sn:0 {0}(952,284)(906,284)(906,280){1}
wire w23;    //: /sn:0 {0}(275,-28)(275,17)(355,17){1}
wire w10;    //: /sn:0 {0}(389,77)(389,116)(449,116){1}
wire w54;    //: /sn:0 {0}(952,374)(517,374)(517,343){1}
wire w24;    //: /sn:0 {0}(294,-28)(294,7)(355,7){1}
wire w21;    //: /sn:0 {0}(168,-4)(130,-4)(130,-28){1}
wire w31;    //: /sn:0 {0}(521,-28)(521,18)(588,18){1}
wire [3:0] w1;    //: /sn:0 {0}(275,188)(275,118)(167,118){1}
wire w32;    //: /sn:0 {0}(536,-28)(536,8)(588,8){1}
wire w53;    //: /sn:0 {0}(952,384)(495,384)(495,343){1}
wire [3:0] w46;    //: /sn:0 /dp:1 {0}(800,107)(806,107)(806,190){1}
wire w8;    //: /sn:0 {0}(161,113)(125,113)(125,77){1}
wire w52;    //: /sn:0 {0}(952,394)(481,394)(481,343){1}
wire [3:0] w17;    //: /sn:0 /dp:1 {0}(802,2)(854,2)(854,190){1}
wire w44;    //: /sn:0 {0}(796,-13)(783,-13)(783,-28){1}
wire w27;    //: /sn:0 {0}(355,-13)(331,-13)(331,-28){1}
wire [3:0] w33;    //: /sn:0 /dp:1 {0}(594,3)(689,3)(689,192){1}
wire w35;    //: /sn:0 {0}(588,-12)(570,-12)(570,-28){1}
wire w28;    //: /sn:0 {0}(687,238)(687,265)(448,265)(448,234){1}
wire w45;    //: /sn:0 {0}(743,77)(743,112)(794,112){1}
wire w14;    //: /sn:0 {0}(725,77)(725,122)(794,122){1}
wire w48;    //: /sn:0 {0}(794,92)(778,92)(778,77){1}
wire w2;    //: /sn:0 {0}(730,-28)(730,17)(796,17){1}
wire w41;    //: /sn:0 {0}(852,236)(852,270)(638,270)(638,238){1}
wire [3:0] w11;    //: /sn:0 /dp:1 {0}(455,111)(468,111)(468,161)(451,161)(451,188){1}
wire w47;    //: /sn:0 {0}(794,102)(761,102)(761,77){1}
wire w15;    //: /sn:0 {0}(99,-28)(99,16)(168,16){1}
wire w61;    //: /sn:0 {0}(952,304)(869,304)(869,280){1}
wire w55;    //: /sn:0 {0}(952,364)(545,364)(545,342){1}
wire w38;    //: /sn:0 {0}(612,105)(580,105)(580,77){1}
wire w5;    //: /sn:0 {0}(84,77)(84,133)(161,133){1}
wire [3:0] w43;    //: /sn:0 {0}(936,276)(906,276){1}
//: {2}(905,276)(887,276){3}
//: {4}(886,276)(869,276){5}
//: {6}(868,276)(839,276){7}
//: {8}(838,276)(831,276)(831,236){9}
wire w26;    //: /sn:0 {0}(355,-3)(314,-3)(314,-28){1}
wire w9;    //: /sn:0 {0}(161,103)(144,103)(144,77){1}
wire w57;    //: /sn:0 {0}(952,344)(692,344)(692,319){1}
wire w51;    //: /sn:0 {0}(952,404)(371,404)(371,377){1}
wire w40;    //: /sn:0 {0}(314,377)(314,434)(952,434){1}
//: enddecls

  tran g44(.Z(w47), .I(A[14]));   //: @(761,71) /sn:0 /R:1 /w:[ 1 29 30 ] /ss:1
  tran g8(.Z(w5), .I(A[0]));   //: @(84,71) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  concat g4 (.I0(w5), .I1(w6), .I2(w8), .I3(w9), .Z(w1));   //: @(166,118) /sn:0 /w:[ 1 1 0 0 1 ] /dr:0
  //: output g47 (Cout) @(928,261) /sn:0 /w:[ 1 ]
  tran g16(.Z(w22), .I(B[3]));   //: @(147,-34) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  CPA2 g3 (.A(w1), .B(w20), .Cin(Cin), .S(w4), .Cout(w16));   //: @(259, 189) /sz:(88, 44) /sn:0 /p:[ Ti0>0 Ti1>1 Bi0>0 Bo0<0 Bo1<1 ]
  concat g26 (.I0(w31), .I1(w32), .I2(w34), .I3(w35), .Z(w33));   //: @(593,3) /sn:0 /w:[ 1 1 0 0 0 ] /dr:0
  tran g17(.Z(w21), .I(B[2]));   //: @(130,-34) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g2 (Cin) @(178,281) /sn:0 /w:[ 1 ]
  tran g30(.Z(w31), .I(B[8]));   //: @(521,-34) /sn:0 /R:1 /w:[ 0 17 18 ] /ss:1
  tran g23(.Z(w24), .I(B[5]));   //: @(294,-34) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1
  tran g39(.Z(w29), .I(B[14]));   //: @(763,-34) /sn:0 /R:1 /w:[ 1 29 30 ] /ss:1
  tran g24(.Z(w23), .I(B[4]));   //: @(275,-34) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  //: input g1 (B) @(37,-32) /sn:0 /w:[ 0 ]
  tran g60(.Z(w58), .I(w30[2]));   //: @(714,313) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g29(.Z(w32), .I(B[9]));   //: @(536,-34) /sn:0 /R:1 /w:[ 0 19 20 ] /ss:1
  tran g51(.Z(w50), .I(w4[2]));   //: @(353,371) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g18(.Z(w19), .I(B[1]));   //: @(112,-34) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g65(.Z(w63), .I(w43[3]));   //: @(906,274) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  CPA2 g25 (.A(w37), .B(w33), .Cin(w28), .S(w30), .Cout(w41));   //: @(625, 193) /sz:(88, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Bi0>0 Bo0<0 Bo1<1 ]
  tran g10(.Z(w13), .I(A[7]));   //: @(425,71) /sn:0 /R:1 /w:[ 1 15 16 ] /ss:1
  tran g64(.Z(w62), .I(w43[2]));   //: @(887,274) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  concat g49 (.I0(w40), .I1(w42), .I2(w50), .I3(w51), .I4(w52), .I5(w53), .I6(w54), .I7(w55), .I8(w56), .I9(w57), .I10(w58), .I11(w59), .I12(w60), .I13(w61), .I14(w62), .I15(w63), .Z(S));   //: @(957,359) /sn:0 /w:[ 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /dr:0
  tran g50(.Z(w51), .I(w4[3]));   //: @(371,371) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g6(.Z(w8), .I(A[2]));   //: @(125,71) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g58(.Z(w56), .I(w30[0]));   //: @(676,313) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g56(.Z(w54), .I(w18[2]));   //: @(517,337) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g35(.Z(w0), .I(A[8]));   //: @(541,71) /sn:0 /R:1 /w:[ 0 17 18 ] /ss:1
  concat g9 (.I0(w7), .I1(w10), .I2(w12), .I3(w13), .Z(w11));   //: @(454,111) /sn:0 /w:[ 1 1 0 0 0 ] /dr:0
  tran g7(.Z(w6), .I(A[1]));   //: @(101,71) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g59(.Z(w57), .I(w30[1]));   //: @(692,313) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  concat g31 (.I0(w0), .I1(w36), .I2(w38), .I3(w39), .Z(w37));   //: @(617,110) /sn:0 /w:[ 1 1 0 0 0 ] /dr:0
  tran g22(.Z(w26), .I(B[6]));   //: @(314,-34) /sn:0 /R:1 /w:[ 1 13 14 ] /ss:1
  tran g54(.Z(w52), .I(w18[0]));   //: @(481,337) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  tran g45(.Z(w45), .I(A[13]));   //: @(743,71) /sn:0 /R:1 /w:[ 0 27 28 ] /ss:1
  tran g41(.Z(w2), .I(B[12]));   //: @(730,-34) /sn:0 /R:1 /w:[ 0 25 26 ] /ss:1
  CPA2 g36 (.A(w46), .B(w17), .Cin(w41), .S(w43), .Cout(Cout));   //: @(790, 191) /sz:(88, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Bi0>0 Bo0<9 Bo1<0 ]
  tran g33(.Z(w38), .I(A[10]));   //: @(580,71) /sn:0 /R:1 /w:[ 1 21 22 ] /ss:1
  tran g52(.Z(w42), .I(w4[1]));   //: @(334,371) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  concat g42 (.I0(w14), .I1(w45), .I2(w47), .I3(w48), .Z(w46));   //: @(799,107) /sn:0 /w:[ 1 1 0 0 0 ] /dr:0
  tran g40(.Z(w3), .I(B[13]));   //: @(747,-34) /sn:0 /R:1 /w:[ 0 27 28 ] /ss:1
  tran g12(.Z(w10), .I(A[5]));   //: @(389,71) /sn:0 /R:1 /anc:1 /w:[ 0 11 12 ] /ss:1
  tran g57(.Z(w55), .I(w18[3]));   //: @(545,336) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g46(.Z(w14), .I(A[12]));   //: @(725,71) /sn:0 /R:1 /w:[ 0 25 26 ] /ss:1
  tran g34(.Z(w36), .I(A[9]));   //: @(558,71) /sn:0 /R:1 /w:[ 0 19 20 ] /ss:1
  tran g28(.Z(w34), .I(B[10]));   //: @(553,-34) /sn:0 /R:1 /w:[ 1 21 22 ] /ss:1
  CPA2 g14 (.A(w11), .B(w25), .Cin(w16), .S(w18), .Cout(w28));   //: @(435, 189) /sz:(88, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Bi0>0 Bo0<9 Bo1<1 ]
  tran g11(.Z(w12), .I(A[6]));   //: @(408,71) /sn:0 /R:1 /w:[ 1 13 14 ] /ss:1
  tran g5(.Z(w9), .I(A[3]));   //: @(144,71) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g61(.Z(w59), .I(w30[3]));   //: @(737,313) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g21(.Z(w27), .I(B[7]));   //: @(331,-34) /sn:0 /R:1 /w:[ 1 15 16 ] /ss:1
  tran g19(.Z(w15), .I(B[0]));   //: @(99,-34) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g32(.Z(w39), .I(A[11]));   //: @(597,71) /sn:0 /R:1 /w:[ 1 23 24 ] /ss:1
  concat g20 (.I0(w23), .I1(w24), .I2(w26), .I3(w27), .Z(w25));   //: @(360,2) /sn:0 /w:[ 1 1 0 0 0 ] /dr:0
  tran g63(.Z(w61), .I(w43[1]));   //: @(869,274) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  tran g43(.Z(w48), .I(A[15]));   //: @(778,71) /sn:0 /R:1 /w:[ 1 31 32 ] /ss:1
  tran g38(.Z(w44), .I(B[15]));   //: @(783,-34) /sn:0 /R:1 /w:[ 1 31 32 ] /ss:1
  concat g15 (.I0(w15), .I1(w19), .I2(w21), .I3(w22), .Z(w20));   //: @(173,1) /sn:0 /w:[ 1 1 0 0 0 ] /dr:0
  //: input g0 (A) @(37,73) /sn:0 /w:[ 0 ]
  //: output g48 (S) @(999,359) /sn:0 /w:[ 1 ]
  tran g27(.Z(w35), .I(B[11]));   //: @(570,-34) /sn:0 /R:1 /w:[ 1 23 24 ] /ss:1
  tran g62(.Z(w60), .I(w43[0]));   //: @(839,274) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  concat g37 (.I0(w2), .I1(w3), .I2(w29), .I3(w44), .Z(w17));   //: @(801,2) /sn:0 /w:[ 1 1 0 0 0 ] /dr:0
  tran g55(.Z(w53), .I(w18[1]));   //: @(495,337) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  tran g53(.Z(w40), .I(w4[0]));   //: @(314,371) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g13(.Z(w7), .I(A[4]));   //: @(368,71) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1

endmodule

module CPA2(S, A, Cin, B, Cout);
//: interface  /sz:(88, 44) /bd:[ Ti0>B[3:0](64/88) Ti1>A[3:0](16/88) Bi0>Cin(62/88) Bo0<Cout(13/88) Bo1<S[3:0](41/88) ]
input [3:0] B;    //: /sn:0 {0}(-193,252)(-93,252)(-93,261)(-47,261)(-47,245)(-21,245){1}
//: {2}(-20,245)(63,245){3}
//: {4}(64,245)(139,245){5}
//: {6}(140,245)(211,245){7}
//: {8}(212,245)(220,245){9}
input [3:0] A;    //: /sn:0 {0}(-186,168)(-88,168)(-88,192)(-43,192){1}
//: {2}(-42,192)(53,192){3}
//: {4}(54,192)(130,192){5}
//: {6}(131,192)(203,192){7}
//: {8}(204,192)(217,192){9}
input Cin;    //: /sn:0 {0}(-9,94)(18,94)(18,104){1}
output Cout;    //: /sn:0 {0}(330,136)(286,136)(286,140)(260,140){1}
output [3:0] S;    //: /sn:0 {0}(317,59)(399,59)(399,38)(409,38){1}
wire w6;    //: /sn:0 {0}(75,120)(54,120)(54,187){1}
wire w16;    //: /sn:0 {0}(218,121)(204,121)(204,187){1}
wire w7;    //: /sn:0 {0}(75,136)(64,136)(64,240){1}
wire w4;    //: /sn:0 /dp:1 {0}(311,74)(48,74)(48,120)(40,120){1}
wire w20;    //: /sn:0 {0}(311,44)(268,44)(268,123)(260,123){1}
wire w12;    //: /sn:0 {0}(146,138)(140,138)(140,240){1}
wire w19;    //: /sn:0 {0}(311,54)(192,54)(192,124)(188,124){1}
wire w10;    //: /sn:0 {0}(166,108)(166,97)(133,97)(133,139)(117,139){1}
wire w1;    //: /sn:0 {0}(-2,118)(-42,118)(-42,187){1}
wire w17;    //: /sn:0 {0}(218,137)(212,137)(212,240){1}
wire w2;    //: /sn:0 {0}(-2,134)(-20,134)(-20,240){1}
wire w11;    //: /sn:0 {0}(146,122)(131,122)(131,187){1}
wire w15;    //: /sn:0 {0}(238,107)(238,97)(202,97)(202,141)(188,141){1}
wire w5;    //: /sn:0 {0}(95,106)(95,97)(58,97)(58,137)(40,137){1}
wire w9;    //: /sn:0 /dp:1 {0}(311,64)(124,64)(124,122)(117,122){1}
//: enddecls

  FA g4 (.Cin(w5), .B(w7), .A(w6), .Cout(w10), .S(w9));   //: @(76, 107) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Li0>0 Li1>0 Ro0<1 Ro1<1 ]
  tran g8(.Z(w6), .I(A[1]));   //: @(54,190) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:0
  FA g3 (.Cin(Cin), .B(w2), .A(w1), .Cout(w5), .S(w4));   //: @(-1, 105) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Li0>0 Li1>0 Ro0<1 Ro1<1 ]
  //: output g16 (S) @(406,38) /sn:0 /w:[ 1 ]
  concat g17 (.I0(w4), .I1(w9), .I2(w19), .I3(w20), .Z(S));   //: @(316,59) /sn:0 /w:[ 0 0 0 0 0 ] /dr:0
  //: input g2 (A) @(-188,168) /sn:0 /w:[ 0 ]
  //: input g1 (Cin) @(-11,94) /sn:0 /w:[ 0 ]
  tran g10(.Z(w16), .I(A[3]));   //: @(204,190) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:0
  FA g6 (.Cin(w15), .B(w17), .A(w16), .Cout(Cout), .S(w20));   //: @(219, 108) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Li0>0 Li1>0 Ro0<1 Ro1<1 ]
  tran g7(.Z(w1), .I(A[0]));   //: @(-42,190) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:0
  tran g9(.Z(w11), .I(A[2]));   //: @(131,190) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:0
  tran g12(.Z(w2), .I(B[0]));   //: @(-20,243) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:0
  FA g5 (.Cin(w10), .B(w12), .A(w11), .Cout(w15), .S(w19));   //: @(147, 109) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Li0>0 Li1>0 Ro0<1 Ro1<1 ]
  tran g14(.Z(w12), .I(B[2]));   //: @(140,243) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:0
  //: input g11 (B) @(-195,252) /sn:0 /w:[ 0 ]
  //: output g0 (Cout) @(327,136) /sn:0 /w:[ 0 ]
  tran g15(.Z(w17), .I(B[3]));   //: @(212,243) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:0
  tran g13(.Z(w7), .I(B[1]));   //: @(64,243) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:0

endmodule

module main;    //: root_module
wire w4;    //: /sn:0 {0}(206,212)(269,212)(269,209)(279,209){1}
wire [15:0] w0;    //: /sn:0 /dp:1 {0}(432,54)(432,157)(378,157)(378,167){1}
wire w3;    //: /sn:0 {0}(326,239)(326,275){1}
wire [15:0] w1;    //: /sn:0 {0}(548,282)(375,282)(375,239){1}
wire [15:0] w5;    //: /sn:0 /dp:1 {0}(136,88)(136,146)(312,146)(312,167){1}
//: enddecls

  //: switch g4 (w4) @(189,212) /sn:0 /w:[ 0 ] /st:1
  led g3 (.I(w1));   //: @(555,282) /sn:0 /R:3 /w:[ 0 ] /type:2
  //: dip g2 (w0) @(432,44) /sn:0 /w:[ 0 ] /st:22
  //: dip g1 (w5) @(136,78) /sn:0 /w:[ 0 ] /st:36
  led g5 (.I(w3));   //: @(326,282) /sn:0 /R:2 /w:[ 1 ] /type:0
  CPA16 g0 (.B(w0), .A(w5), .Cin(w4), .S(w1), .Cout(w3));   //: @(280, 168) /sz:(144, 70) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Bo1<0 ]

endmodule

module FA(Cout, S, Cin, B, A);
//: interface  /sz:(40, 40) /bd:[ Ti0>Cin(19/40) Li0>B(29/40) Li1>A(13/40) Ro0<Cout(32/40) Ro1<S(15/40) ]
input B;    //: /sn:0 {0}(160,154)(128,154)(128,104)(115,104){1}
//: {2}(113,102)(113,91)(123,91){3}
//: {4}(111,104)(95,104){5}
input A;    //: /sn:0 {0}(97,85)(102,85){1}
//: {2}(106,85)(113,85)(113,86)(123,86){3}
//: {4}(104,87)(104,159)(160,159){5}
input Cin;    //: /sn:0 {0}(99,123)(154,123){1}
//: {2}(156,121)(156,100)(170,100){3}
//: {4}(156,125)(156,129)(160,129){5}
output Cout;    //: /sn:0 {0}(277,142)(233,142){1}
output S;    //: /sn:0 {0}(275,100)(201,100)(201,98)(191,98){1}
wire w13;    //: /sn:0 /dp:1 {0}(212,144)(191,144)(191,157)(181,157){1}
wire w7;    //: /sn:0 {0}(160,134)(149,134)(149,91){1}
//: {2}(151,89)(153,89)(153,95)(170,95){3}
//: {4}(147,89)(144,89){5}
wire w12;    //: /sn:0 /dp:1 {0}(212,139)(191,139)(191,132)(181,132){1}
//: enddecls

  //: output g4 (Cout) @(274,142) /sn:0 /w:[ 0 ]
  and g8 (.I0(B), .I1(A), .Z(w13));   //: @(171,157) /sn:0 /w:[ 0 5 1 ]
  //: output g3 (S) @(272,100) /sn:0 /w:[ 0 ]
  //: input g2 (Cin) @(97,123) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(93,104) /sn:0 /w:[ 5 ]
  //: joint g10 (Cin) @(156, 123) /w:[ -1 2 1 4 ]
  xor g6 (.I0(w7), .I1(Cin), .Z(S));   //: @(181,98) /sn:0 /w:[ 3 3 1 ]
  and g7 (.I0(Cin), .I1(w7), .Z(w12));   //: @(171,132) /sn:0 /w:[ 5 0 1 ]
  or g9 (.I0(w12), .I1(w13), .Z(Cout));   //: @(223,142) /sn:0 /w:[ 0 0 1 ]
  //: joint g12 (A) @(104, 85) /w:[ 2 -1 1 4 ]
  xor g5 (.I0(A), .I1(B), .Z(w7));   //: @(134,89) /sn:0 /w:[ 3 3 5 ]
  //: joint g11 (w7) @(149, 89) /w:[ 2 -1 4 1 ]
  //: input g0 (A) @(95,85) /sn:0 /w:[ 0 ]
  //: joint g13 (B) @(113, 104) /w:[ 1 2 4 -1 ]

endmodule
