//: version "1.8.7"

module FA2(B, A, Cin, Cout, S);
//: interface  /sz:(40, 40) /bd:[ Li0>Cin(7/40) Li1>B(23/40) Li2>A(34/40) Ro0<Cout(31/40) Ro1<S(13/40) ]
input B;    //: /sn:0 {0}(82,83)(73,83)(73,91)(-46,91)(-46,61){1}
//: {2}(-44,59)(-39,59)(-39,35)(6,35){3}
//: {4}(-48,59)(-52,59){5}
input A;    //: /sn:0 {0}(-46,9)(-13,9){1}
//: {2}(-9,9)(-2,9)(-2,30)(6,30){3}
//: {4}(-11,7)(-11,1)(88,1){5}
input Cin;    //: /sn:0 {0}(-55,130)(206,130)(206,123){1}
//: {2}(208,121)(277,121){3}
//: {4}(206,119)(206,90)(219,90){5}
output Cout;    //: /sn:0 {0}(294,178)(410,178){1}
output S;    //: /sn:0 {0}(352,80)(390,80)(390,72)(410,72){1}
wire w4;    //: /sn:0 {0}(166,41)(196,41){1}
//: {2}(200,41)(281,41){3}
//: {4}(198,43)(198,85)(219,85){5}
wire w0;    //: /sn:0 {0}(273,175)(260,175)(260,119){1}
//: {2}(262,117)(268,117)(268,116)(277,116){3}
//: {4}(260,115)(260,90){5}
//: {6}(260,86)(260,46)(281,46){7}
//: {8}(258,88)(240,88){9}
wire w12;    //: /sn:0 {0}(298,119)(320,119)(320,82)(331,82){1}
wire w1;    //: /sn:0 /dp:1 {0}(273,180)(64,180)(64,80){1}
//: {2}(66,78)(82,78){3}
//: {4}(64,76)(64,34){5}
//: {6}(64,30)(64,6)(88,6){7}
//: {8}(62,32)(52,32)(52,33)(27,33){9}
wire w8;    //: /sn:0 {0}(103,81)(135,81)(135,43)(145,43){1}
wire w2;    //: /sn:0 {0}(109,4)(136,4)(136,38)(145,38){1}
wire w5;    //: /sn:0 {0}(302,44)(321,44)(321,77)(331,77){1}
//: enddecls

  //: joint g4 (w1) @(64, 32) /w:[ -1 6 8 5 ]
  nand g8 (.I0(w4), .I1(Cin), .Z(w0));   //: @(230,88) /sn:0 /delay:" 3" /w:[ 5 5 9 ]
  nand g16 (.I0(w0), .I1(w1), .Z(Cout));   //: @(284,178) /sn:0 /delay:" 3" /w:[ 0 0 0 ]
  //: joint g3 (A) @(-11, 9) /w:[ 2 4 1 -1 ]
  //: joint g17 (Cin) @(206, 121) /w:[ 2 4 -1 1 ]
  nand g2 (.I0(w1), .I1(B), .Z(w8));   //: @(93,81) /sn:0 /delay:" 3" /w:[ 3 0 0 ]
  nand g1 (.I0(A), .I1(B), .Z(w1));   //: @(17,33) /sn:0 /delay:" 3" /w:[ 3 3 9 ]
  //: joint g18 (w1) @(64, 78) /w:[ 2 4 -1 1 ]
  //: input g10 (B) @(-54,59) /sn:0 /w:[ 5 ]
  nand g6 (.I0(w2), .I1(w8), .Z(w4));   //: @(156,41) /sn:0 /delay:" 3" /w:[ 1 1 0 ]
  nand g7 (.I0(w4), .I1(w0), .Z(w5));   //: @(292,44) /sn:0 /delay:" 3" /w:[ 3 7 0 ]
  //: input g9 (A) @(-48,9) /sn:0 /w:[ 0 ]
  nand g12 (.I0(w0), .I1(Cin), .Z(w12));   //: @(288,119) /sn:0 /delay:" 3" /w:[ 3 3 0 ]
  //: joint g14 (w0) @(260, 88) /w:[ -1 6 8 5 ]
  //: joint g5 (B) @(-46, 59) /w:[ 2 -1 4 1 ]
  //: input g11 (Cin) @(-57,130) /sn:0 /w:[ 0 ]
  nand g19 (.I0(w5), .I1(w12), .Z(S));   //: @(342,80) /sn:0 /delay:" 3" /w:[ 1 1 0 ]
  //: output g21 (Cout) @(407,178) /sn:0 /w:[ 1 ]
  //: output g20 (S) @(407,72) /sn:0 /w:[ 1 ]
  //: joint g15 (w0) @(260, 117) /w:[ 2 4 -1 1 ]
  nand g0 (.I0(A), .I1(w1), .Z(w2));   //: @(99,4) /sn:0 /delay:" 3" /w:[ 5 7 0 ]
  //: joint g13 (w4) @(198, 41) /w:[ 2 -1 1 4 ]

endmodule

module main;    //: root_module
wire w4;    //: /sn:0 {0}(395,281)(435,281)(435,312)(445,312){1}
wire w0;    //: /sn:0 {0}(131,183)(262,183)(262,237)(272,237){1}
wire w3;    //: /sn:0 {0}(395,248)(446,248)(446,198){1}
wire w1;    //: /sn:0 /dp:1 {0}(272,266)(157,266){1}
wire w5;    //: /sn:0 {0}(111,348)(262,348)(262,287)(272,287){1}
//: enddecls

  led g4 (.I(w3));   //: @(446,191) /sn:0 /w:[ 1 ] /type:0
  //: switch g3 (w0) @(114,183) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w1) @(140,266) /sn:0 /w:[ 1 ] /st:0
  FA2 g1 (.Cin(w0), .B(w1), .A(w5), .Cout(w4), .S(w3));   //: @(273, 225) /sz:(121, 73) /sn:0 /p:[ Li0>1 Li1>0 Li2>1 Ro0<0 Ro1<0 ]
  led g5 (.I(w4));   //: @(452,312) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: switch g0 (w5) @(94,348) /sn:0 /w:[ 0 ] /st:0

endmodule
