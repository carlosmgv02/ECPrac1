//: version "1.8.7"

module FullAdder(A, Cin, B, S, Cout);
//: interface  /sz:(96, 73) /bd:[ Ti0>A(22/96) Ti1>B(63/96) Li0>Cin(30/73) Bo0<S(31/96) Bo1<Cout(61/96) ]
input B;    //: /sn:0 {0}(93,188)(27,188)(27,124){1}
//: {2}(29,122)(35,122){3}
//: {4}(25,122)(9,122)(9,125)(-12,125){5}
input A;    //: /sn:0 {0}(-12,110)(8,110)(8,117)(14,117){1}
//: {2}(18,117)(35,117){3}
//: {4}(16,119)(16,193)(93,193){5}
input Cin;    //: /sn:0 {0}(-13,143)(80,143){1}
//: {2}(82,141)(82,125)(91,125){3}
//: {4}(82,145)(82,163)(92,163){5}
output Cout;    //: /sn:0 {0}(165,179)(193,179){1}
output S;    //: /sn:0 {0}(112,123)(167,123){1}
wire w14;    //: /sn:0 {0}(56,120)(63,120){1}
//: {2}(67,120)(91,120){3}
//: {4}(65,122)(65,168)(92,168){5}
wire w2;    //: /sn:0 {0}(114,191)(134,191)(134,181)(144,181){1}
wire w5;    //: /sn:0 {0}(113,166)(134,166)(134,176)(144,176){1}
//: enddecls

  //: input g8 (A) @(-14,110) /sn:0 /w:[ 0 ]
  xor g4 (.I0(A), .I1(B), .Z(w14));   //: @(46,120) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  xor g3 (.I0(w14), .I1(Cin), .Z(S));   //: @(102,123) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  or g2 (.I0(w5), .I1(w2), .Z(Cout));   //: @(155,179) /sn:0 /w:[ 1 1 0 ]
  and g1 (.I0(Cin), .I1(w14), .Z(w5));   //: @(103,166) /sn:0 /delay:" 1" /w:[ 5 5 0 ]
  //: input g10 (Cin) @(-15,143) /sn:0 /w:[ 0 ]
  //: joint g6 (B) @(27, 122) /w:[ 2 -1 4 1 ]
  //: input g9 (B) @(-14,125) /sn:0 /w:[ 5 ]
  //: joint g7 (A) @(16, 117) /w:[ 2 -1 1 4 ]
  //: output g12 (S) @(164,123) /sn:0 /w:[ 1 ]
  //: joint g11 (Cin) @(82, 143) /w:[ -1 2 1 4 ]
  //: joint g5 (w14) @(65, 120) /w:[ 2 -1 1 4 ]
  and g0 (.I0(B), .I1(A), .Z(w2));   //: @(104,191) /sn:0 /w:[ 0 5 0 ]
  //: output g13 (Cout) @(190,179) /sn:0 /w:[ 1 ]

endmodule

module main;    //: root_module
wire w3;    //: /sn:0 {0}(194,249)(194,228){1}
wire w0;    //: /sn:0 {0}(182,98)(196,98)(196,153){1}
wire w10;    //: /sn:0 {0}(135,120)(155,120)(155,153){1}
wire w1;    //: /sn:0 {0}(111,184)(132,184){1}
wire w2;    //: /sn:0 {0}(164,248)(164,228){1}
wire w11;    //: /sn:0 {0}(-28251,189)(-28251,199){1}
//: enddecls

  //: switch g4 (w0) @(165,98) /sn:0 /w:[ 0 ] /st:1
  //: switch g3 (w11) @(-28251,176) /sn:0 /R:3 /w:[ 0 ] /st:0
  //: switch g2 (w10) @(118,120) /sn:0 /w:[ 0 ] /st:1
  led g1 (.I(w2));   //: @(164,255) /sn:0 /R:2 /w:[ 0 ] /type:0
  led g6 (.I(w3));   //: @(194,256) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: switch g5 (w1) @(94,184) /sn:0 /w:[ 0 ] /st:0
  FullAdder g0 (.B(w0), .A(w10), .Cin(w1), .Cout(w3), .S(w2));   //: @(133, 154) /sz:(96, 73) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Bo1<1 ]

endmodule
