//: version "1.8.7"

module HA(CO, S, B, A);
//: interface  /sz:(133, 96) /bd:[ Ti0>A(39/133) Bi0>B(39/133) Ro0<CO(43/96) Ro1<S(60/96) ]
input B;    //: /sn:0 /dp:1 {0}(287,136)(248,136)(248,156)(215,156){1}
//: {2}(211,156)(178,156)(178,211)(175,211){3}
//: {4}(213,158)(213,218)(278,218)(278,212)(288,212){5}
input A;    //: /sn:0 {0}(186,129)(203,129)(203,126)(225,126){1}
//: {2}(229,126)(274,126)(274,131)(287,131){3}
//: {4}(227,128)(227,207)(288,207){5}
output CO;    //: /sn:0 /dp:1 {0}(309,210)(412,210)(412,216)(422,216){1}
output S;    //: /sn:0 /dp:1 {0}(308,134)(418,134)(418,122)(428,122){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(298,134) /sn:0 /w:[ 3 0 0 ]
  //: output g3 (CO) @(419,216) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(425,122) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(173,211) /sn:0 /w:[ 3 ]
  //: joint g6 (B) @(213, 156) /w:[ 1 -1 2 4 ]
  //: joint g7 (A) @(227, 126) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(CO));   //: @(299,210) /sn:0 /w:[ 5 5 0 ]
  //: input g0 (A) @(184,129) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire w0;    //: /sn:0 {0}(454,220)(454,230)(408,230){1}
wire w3;    //: /sn:0 {0}(263,339)(313,339)(313,284){1}
wire w1;    //: /sn:0 {0}(446,252)(446,266)(424,266)(424,247)(408,247){1}
wire w2;    //: /sn:0 {0}(302,150)(313,150)(313,186){1}
//: enddecls

  //: switch g4 (w3) @(246,339) /sn:0 /w:[ 0 ] /st:1
  //: switch g3 (w2) @(285,150) /sn:0 /w:[ 0 ] /st:0
  led g2 (.I(w1));   //: @(446,245) /sn:0 /w:[ 0 ] /type:0
  led g1 (.I(w0));   //: @(454,213) /sn:0 /w:[ 0 ] /type:0
  HA g0 (.A(w2), .B(w3), .CO(w0), .S(w1));   //: @(274, 187) /sz:(133, 96) /sn:0 /p:[ Ti0>1 Bi0>1 Ro0<1 Ro1<1 ]

endmodule
