//: version "1.8.7"

module PFA(Pi, S, Ci, B, Gi, A);
//: interface  /sz:(40, 40) /bd:[ Li0>Ci(37/40) Li1>B(23/40) Li2>A(8/40) Ro0<Gi(37/40) Ro1<Pi(26/40) Ro2<S(12/40) ]
input B;    //: /sn:0 {0}(206,145)(223,145){1}
//: {2}(227,145)(269,145)(269,133)(279,133){3}
//: {4}(225,147)(225,188){5}
//: {6}(227,190)(354,190){7}
//: {8}(225,192)(225,229)(356,229){9}
output Gi;    //: /sn:0 {0}(435,225)(387,225)(387,227)(377,227){1}
input A;    //: /sn:0 {0}(205,117)(246,117){1}
//: {2}(250,117)(269,117)(269,128)(279,128){3}
//: {4}(248,119)(248,183){5}
//: {6}(250,185)(354,185){7}
//: {8}(248,187)(248,224)(356,224){9}
output Pi;    //: /sn:0 /dp:1 {0}(375,188)(422,188)(422,187)(432,187){1}
input Ci;    //: /sn:0 /dp:1 {0}(351,146)(314,146)(314,174)(204,174){1}
output S;    //: /sn:0 /dp:1 {0}(372,144)(423,144)(423,145)(433,145){1}
wire w2;    //: /sn:0 {0}(300,131)(341,131)(341,141)(351,141){1}
//: enddecls

  //: output g4 (Pi) @(429,187) /sn:0 /w:[ 1 ]
  or g8 (.I0(A), .I1(B), .Z(Pi));   //: @(365,188) /sn:0 /delay:" 3" /w:[ 7 7 0 ]
  //: output g3 (S) @(430,145) /sn:0 /w:[ 1 ]
  //: input g2 (Ci) @(202,174) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(204,145) /sn:0 /w:[ 0 ]
  //: joint g10 (A) @(248, 117) /w:[ 2 -1 1 4 ]
  xor g6 (.I0(A), .I1(B), .Z(w2));   //: @(290,131) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  xor g7 (.I0(w2), .I1(Ci), .Z(S));   //: @(362,144) /sn:0 /delay:" 4" /w:[ 1 0 0 ]
  and g9 (.I0(A), .I1(B), .Z(Gi));   //: @(367,227) /sn:0 /delay:" 3" /w:[ 9 9 1 ]
  //: joint g12 (B) @(225, 145) /w:[ 2 -1 1 4 ]
  //: output g5 (Gi) @(432,225) /sn:0 /w:[ 0 ]
  //: joint g11 (A) @(248, 185) /w:[ 6 5 -1 8 ]
  //: input g0 (A) @(203,117) /sn:0 /w:[ 0 ]
  //: joint g13 (B) @(225, 190) /w:[ 6 5 -1 8 ]

endmodule

module main;    //: root_module
wire w4;    //: /sn:0 /dp:1 {0}(404,168)(404,185)(328,185){1}
wire w3;    //: /sn:0 /dp:1 {0}(389,99)(389,165)(328,165){1}
wire w0;    //: /sn:0 {0}(91,155)(250,155)(250,180)(270,180){1}
wire w1;    //: /sn:0 {0}(110,208)(250,208)(250,198)(270,198){1}
wire w8;    //: /sn:0 {0}(270,159)(251,159)(251,149)(241,149)(241,97)(159,97){1}
wire w5;    //: /sn:0 /dp:1 {0}(413,211)(408,211)(408,198)(328,198){1}
//: enddecls

  //: switch g4 (w0) @(74,155) /sn:0 /w:[ 0 ] /st:0
  //: switch g3 (w8) @(142,97) /sn:0 /w:[ 1 ] /st:0
  led g2 (.I(w5));   //: @(420,211) /sn:0 /R:3 /w:[ 0 ] /type:0
  led g1 (.I(w4));   //: @(404,161) /sn:0 /w:[ 0 ] /type:0
  led g6 (.I(w3));   //: @(389,92) /sn:0 /w:[ 0 ] /type:0
  //: switch g5 (w1) @(93,208) /sn:0 /w:[ 0 ] /st:0
  PFA g0 (.A(w8), .B(w0), .Ci(w1), .S(w3), .Pi(w4), .Gi(w5));   //: @(271, 149) /sz:(56, 54) /sn:0 /p:[ Li0>0 Li1>1 Li2>1 Ro0<1 Ro1<1 Ro2<1 ]

endmodule
