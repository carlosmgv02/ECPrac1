//: version "1.8.7"

module CLA_2(S, GG, A, B, C0, PG);
//: interface  /sz:(99, 96) /bd:[ Ti0>B[3:0](71/99) Ti1>A[3:0](13/99) Li0>C0(49/96) Bo0<S(83/99) Bo1<GG(49/99) Bo2<PG(24/99) ]
input [3:0] B;    //: /sn:0 {0}(937,92)(834,92){1}
//: {2}(833,92)(652,92){3}
//: {4}(651,92)(491,92){5}
//: {6}(490,92)(315,92){7}
//: {8}(314,92)(116,92){9}
input C0;    //: /sn:0 {0}(224,226)(236,226){1}
//: {2}(240,226)(259,226)(259,225)(267,225){3}
//: {4}(238,228)(238,374)(259,374){5}
output GG;    //: /sn:0 {0}(1014,390)(899,390){1}
input [3:0] A;    //: /sn:0 {0}(121,67)(276,67){1}
//: {2}(277,67)(458,67){3}
//: {4}(459,67)(537,67)(537,66)(616,66){5}
//: {6}(617,66)(785,66){7}
//: {8}(786,66)(931,66){9}
output PG;    //: /sn:0 {0}(1012,366)(899,366){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(986,545)(1031,545){1}
wire w6;    //: /sn:0 {0}(459,179)(459,71){1}
wire w13;    //: /sn:0 {0}(664,178)(664,104)(652,104)(652,96){1}
wire w7;    //: /sn:0 {0}(495,179)(495,104)(491,104)(491,96){1}
wire w34;    //: /sn:0 /dp:1 {0}(414,348)(414,226)(444,226){1}
wire w0;    //: /sn:0 {0}(282,178)(282,79)(277,79)(277,71){1}
wire w3;    //: /sn:0 {0}(329,277)(329,305)(306,305)(306,320)(300,320)(300,348){1}
wire w22;    //: /sn:0 {0}(885,210)(919,210)(919,530)(980,530){1}
wire w30;    //: /sn:0 /dp:1 {0}(648,348)(648,287)(675,287)(675,277){1}
wire w12;    //: /sn:0 {0}(628,178)(628,78)(617,78)(617,70){1}
wire w18;    //: /sn:0 {0}(798,177)(798,78)(786,78)(786,70){1}
wire w19;    //: /sn:0 {0}(834,177)(834,96){1}
wire w23;    //: /sn:0 {0}(885,245)(895,245)(895,305)(850,305)(850,348){1}
wire w1;    //: /sn:0 {0}(318,178)(318,104)(315,104)(315,96){1}
wire w31;    //: /sn:0 /dp:1 {0}(592,348)(592,225)(613,225){1}
wire w32;    //: /sn:0 /dp:1 {0}(504,348)(504,326)(561,326)(561,247)(546,247){1}
wire w8;    //: /sn:0 /dp:1 {0}(980,550)(576,550)(576,212)(546,212){1}
wire w17;    //: /sn:0 {0}(715,246)(731,246)(731,330)(690,330)(690,348){1}
wire w27;    //: /sn:0 /dp:1 {0}(825,348)(825,286)(845,286)(845,276){1}
wire w28;    //: /sn:0 /dp:1 {0}(767,348)(767,224)(783,224){1}
wire w33;    //: /sn:0 /dp:1 {0}(464,348)(464,288)(506,288)(506,278){1}
wire w2;    //: /sn:0 /dp:1 {0}(980,560)(387,560)(387,211)(369,211){1}
wire w11;    //: /sn:0 {0}(980,540)(748,540)(748,211)(715,211){1}
wire w5;    //: /sn:0 {0}(369,246)(392,246)(392,295)(342,295)(342,320)(329,320)(329,348){1}
//: enddecls

  CLL_2 g4 (.G0(w3), .P0(w5), .G1(w33), .P1(w32), .G2(w30), .P2(w17), .G3(w27), .P3(w23), .C0(C0), .C1(w34), .C2(w31), .C3(w28), .GG(GG), .PG(PG));   //: @(260, 349) /sz:(638, 57) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>0 Ti3>0 Ti4>0 Ti5>1 Ti6>0 Ti7>1 Li0>5 To0<0 To1<0 To2<0 Ro0<1 Ro1<1 ]
  tran g8(.Z(w0), .I(A[0]));   //: @(277,65) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  PFA g3 (.B(w19), .A(w18), .Ci(w28), .Gi(w27), .Pi(w23), .S(w22));   //: @(784, 178) /sz:(100, 97) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<0 Ro1<0 ]
  //: joint g16 (C0) @(238, 226) /w:[ 2 -1 1 4 ]
  //: output g17 (S) @(1028,545) /sn:0 /w:[ 1 ]
  PFA g2 (.B(w13), .A(w12), .Ci(w31), .Gi(w30), .Pi(w17), .S(w11));   //: @(614, 179) /sz:(100, 97) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<0 Ro1<1 ]
  PFA g1 (.B(w7), .A(w6), .Ci(w34), .Gi(w33), .Pi(w32), .S(w8));   //: @(445, 180) /sz:(100, 97) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<1 Ro1<1 ]
  //: output g18 (GG) @(1011,390) /sn:0 /w:[ 0 ]
  tran g10(.Z(w6), .I(A[1]));   //: @(459,65) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: input g6 (A) @(119,67) /sn:0 /w:[ 0 ]
  //: input g7 (B) @(114,92) /sn:0 /w:[ 9 ]
  tran g9(.Z(w1), .I(B[0]));   //: @(315,90) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  tran g12(.Z(w12), .I(A[2]));   //: @(617,64) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g5 (C0) @(222,226) /sn:0 /w:[ 0 ]
  tran g11(.Z(w7), .I(B[1]));   //: @(491,90) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  tran g14(.Z(w18), .I(A[3]));   //: @(786,64) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: output g19 (PG) @(1009,366) /sn:0 /w:[ 0 ]
  concat g20 (.I0(w2), .I1(w8), .I2(w11), .I3(w22), .Z(S));   //: @(985,545) /sn:0 /w:[ 0 0 0 1 0 ] /dr:0
  PFA g0 (.B(w1), .A(w0), .Ci(C0), .Gi(w3), .Pi(w5), .S(w2));   //: @(268, 179) /sz:(100, 97) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>3 Bo0<0 Ro0<0 Ro1<1 ]
  tran g15(.Z(w19), .I(B[3]));   //: @(834,90) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g13(.Z(w13), .I(B[2]));   //: @(652,90) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1

endmodule

module CLU_16(P2, C0, P1, GG, G1, C1, G0, C2, C3, C4, P3, G3, PG, G2, P0);
//: interface  /sz:(40, 40) /bd:[ ]
input G2;    //: /sn:0 {0}(361,21)(340,21)(340,64)(-38,64){1}
//: {2}(-40,62)(-40,-203){3}
//: {4}(-40,66)(-40,248)(229,248){5}
input C0;    //: /sn:0 /dp:11 {0}(249,-29)(191,-29)(191,-39)(156,-39){1}
//: {2}(154,-41)(154,-126){3}
//: {4}(156,-128)(190,-128)(190,-117)(241,-117){5}
//: {6}(154,-130)(154,-180){7}
//: {8}(156,-182)(195,-182)(195,-189)(242,-189){9}
//: {10}(154,-184)(154,-205){11}
//: {12}(154,-37)(154,101)(225,101){13}
output GG;    //: /sn:0 {0}(389,187)(426,187)(426,201)(436,201){1}
input P1;    //: /sn:0 {0}(225,111)(5,111){1}
//: {2}(3,109)(3,11){3}
//: {4}(5,9)(138,9)(138,10)(247,10){5}
//: {6}(3,7)(3,-21){7}
//: {8}(5,-23)(40,-23)(40,-19)(249,-19){9}
//: {10}(3,-25)(3,-85){11}
//: {12}(5,-87)(40,-87)(40,-84)(242,-84){13}
//: {14}(3,-89)(3,-106){15}
//: {16}(5,-108)(135,-108)(135,-107)(241,-107){17}
//: {18}(3,-110)(3,-209){19}
//: {20}(3,113)(3,146){21}
//: {22}(5,148)(115,148)(115,151)(226,151){23}
//: {24}(3,150)(3,183)(228,183){25}
output C3;    //: /sn:0 {0}(382,13)(426,13)(426,16)(436,16){1}
output PG;    //: /sn:0 {0}(247,153)(420,153)(420,151)(435,151){1}
input G0;    //: /sn:0 {0}(100,-206)(100,-169){1}
//: {2}(102,-167)(174,-167)(174,-168)(362,-168){3}
//: {4}(100,-165)(100,-94){5}
//: {6}(102,-92)(193,-92)(193,-89)(242,-89){7}
//: {8}(100,-90)(100,0){9}
//: {10}(102,2)(196,2)(196,5)(247,5){11}
//: {12}(100,4)(100,178)(228,178){13}
output C4;    //: /sn:0 {0}(389,107)(418,107)(418,109)(433,109){1}
output C2;    //: /sn:0 {0}(378,-87)(426,-87)(426,-85)(436,-85){1}
input P3;    //: /sn:0 {0}(225,121)(48,121)(48,120)(-101,120){1}
//: {2}(-103,118)(-103,-204){3}
//: {4}(-103,122)(-103,157){5}
//: {6}(-101,159)(46,159)(46,161)(226,161){7}
//: {8}(-103,161)(-103,184){9}
//: {10}(-101,186)(-93,186)(-93,193)(228,193){11}
//: {12}(-103,188)(-103,215){13}
//: {14}(-101,217)(-92,217)(-92,223)(229,223){15}
//: {16}(-103,219)(-103,253)(229,253){17}
input G1;    //: /sn:0 {0}(357,-82)(220,-82)(220,-81)(29,-81){1}
//: {2}(27,-83)(27,-215){3}
//: {4}(27,-79)(27,34){5}
//: {6}(29,36)(63,36)(63,39)(249,39){7}
//: {8}(27,38)(27,213)(229,213){9}
input G3;    //: /sn:0 {0}(-125,-203)(-125,276)(315,276){1}
//: {2}(319,276)(363,276)(363,195)(368,195){3}
//: {4}(317,274)(317,117)(368,117){5}
input P0;    //: /sn:0 /dp:15 {0}(225,106)(85,106)(85,102)(75,102){1}
//: {2}(73,100)(73,-26){3}
//: {4}(75,-28)(184,-28)(184,-24)(249,-24){5}
//: {6}(73,-30)(73,-112){7}
//: {8}(75,-114)(170,-114)(170,-112)(241,-112){9}
//: {10}(73,-116)(73,-177){11}
//: {12}(75,-179)(181,-179)(181,-184)(242,-184){13}
//: {14}(73,-181)(73,-205){15}
//: {16}(73,104)(73,146)(226,146){17}
output C1;    //: /sn:0 {0}(383,-170)(426,-170)(426,-168)(436,-168){1}
input P2;    //: /sn:0 {0}(225,116)(-51,116)(-51,114)(-61,114){1}
//: {2}(-63,112)(-63,44){3}
//: {4}(-61,42)(106,42)(106,44)(249,44){5}
//: {6}(-63,40)(-63,12){7}
//: {8}(-61,10)(-27,10)(-27,15)(247,15){9}
//: {10}(-63,8)(-63,-15){11}
//: {12}(-61,-17)(97,-17)(97,-14)(249,-14){13}
//: {14}(-63,-19)(-63,-202){15}
//: {16}(-63,116)(-63,153){17}
//: {18}(-61,155)(74,155)(74,156)(226,156){19}
//: {20}(-63,157)(-63,182){21}
//: {22}(-61,184)(-53,184)(-53,188)(228,188){23}
//: {24}(-63,186)(-63,218)(229,218){25}
wire w3;    //: /sn:0 {0}(246,111)(271,111)(271,97)(368,97){1}
wire w23;    //: /sn:0 {0}(249,185)(278,185){1}
//: {2}(282,185)(368,185){3}
//: {4}(280,183)(280,102)(368,102){5}
wire w8;    //: /sn:0 {0}(263,-86)(347,-86)(347,-87)(357,-87){1}
wire G4;    //: /sn:0 {0}(368,112)(301,112)(301,249){1}
//: {2}(303,251)(360,251)(360,190)(368,190){3}
//: {4}(299,251)(250,251){5}
wire w17;    //: /sn:0 {0}(270,42)(327,42)(327,16)(361,16){1}
wire w14;    //: /sn:0 {0}(268,10)(351,10)(351,11)(361,11){1}
wire w11;    //: /sn:0 {0}(270,-22)(351,-22)(351,6)(361,6){1}
wire w2;    //: /sn:0 {0}(263,-186)(342,-186)(342,-173)(362,-173){1}
wire w5;    //: /sn:0 {0}(262,-112)(347,-112)(347,-92)(357,-92){1}
wire w26;    //: /sn:0 {0}(250,218)(290,218){1}
//: {2}(294,218)(340,218)(340,180)(368,180){3}
//: {4}(292,216)(292,107)(368,107){5}
//: enddecls

  //: input g4 (P2) @(-63,-204) /sn:0 /R:3 /w:[ 15 ]
  //: input g8 (C0) @(154,-207) /sn:0 /R:3 /w:[ 11 ]
  //: joint g44 (P2) @(-63, 42) /w:[ 4 6 -1 3 ]
  //: input g3 (P1) @(3,-211) /sn:0 /R:3 /w:[ 19 ]
  and g16 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w23));   //: @(239,185) /sn:0 /w:[ 13 25 23 11 0 ]
  and g17 (.I0(G1), .I1(P2), .I2(P3), .Z(w26));   //: @(240,218) /sn:0 /w:[ 9 25 15 0 ]
  //: output g26 (GG) @(433,201) /sn:0 /w:[ 1 ]
  //: input g2 (G1) @(27,-217) /sn:0 /R:3 /w:[ 3 ]
  //: output g23 (C1) @(433,-168) /sn:0 /w:[ 1 ]
  //: joint g30 (C0) @(154, -128) /w:[ 4 6 -1 3 ]
  //: input g1 (G0) @(100,-208) /sn:0 /R:3 /w:[ 0 ]
  //: joint g39 (P2) @(-63, -17) /w:[ 12 14 -1 11 ]
  //: output g24 (C2) @(433,-85) /sn:0 /w:[ 1 ]
  //: joint g29 (G0) @(100, -167) /w:[ 2 1 -1 4 ]
  //: joint g70 (G4) @(301, 251) /w:[ 2 1 4 -1 ]
  and g18 (.I0(G2), .I1(P3), .Z(G4));   //: @(240,251) /sn:0 /w:[ 5 17 5 ]
  //: joint g65 (P0) @(73, 102) /w:[ 1 2 -1 16 ]
  and g10 (.I0(C0), .I1(P0), .I2(P1), .Z(w5));   //: @(252,-112) /sn:0 /w:[ 5 9 17 0 ]
  //: output g25 (C3) @(433,16) /sn:0 /w:[ 1 ]
  //: joint g64 (P1) @(3, 111) /w:[ 1 2 -1 20 ]
  //: output g72 (C4) @(430,109) /sn:0 /w:[ 1 ]
  //: joint g49 (P2) @(-63, 155) /w:[ 18 17 -1 20 ]
  //: joint g50 (P3) @(-103, 159) /w:[ 6 5 -1 8 ]
  //: input g6 (P3) @(-103,-206) /sn:0 /R:3 /w:[ 3 ]
  //: input g7 (G3) @(-125,-205) /sn:0 /R:3 /w:[ 0 ]
  and g9 (.I0(C0), .I1(P0), .Z(w2));   //: @(253,-186) /sn:0 /w:[ 9 13 0 ]
  //: joint g68 (w23) @(280, 185) /w:[ 2 4 1 -1 ]
  //: joint g35 (G1) @(27, -81) /w:[ 1 2 -1 4 ]
  //: joint g31 (P0) @(73, -114) /w:[ 8 10 -1 7 ]
  //: joint g71 (G3) @(317, 276) /w:[ 2 4 1 -1 ]
  or g22 (.I0(w26), .I1(w23), .I2(G4), .I3(G3), .Z(GG));   //: @(379,187) /sn:0 /w:[ 3 3 3 3 0 ]
  or g67 (.I0(w3), .I1(w23), .I2(w26), .I3(G4), .I4(G3), .Z(C4));   //: @(379,107) /sn:0 /w:[ 1 5 5 0 5 0 ]
  //: joint g36 (C0) @(154, -39) /w:[ 1 2 -1 12 ]
  //: joint g41 (P1) @(3, 9) /w:[ 4 6 -1 3 ]
  //: joint g54 (P3) @(-103, 186) /w:[ 10 9 -1 12 ]
  //: joint g45 (G2) @(-40, 64) /w:[ 1 2 -1 4 ]
  //: joint g33 (G0) @(100, -92) /w:[ 6 5 -1 8 ]
  //: joint g69 (w26) @(292, 218) /w:[ 2 4 1 -1 ]
  //: joint g42 (P2) @(-63, 10) /w:[ 8 10 -1 7 ]
  //: joint g40 (G0) @(100, 2) /w:[ 10 9 -1 12 ]
  and g12 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .Z(w11));   //: @(260,-22) /sn:0 /w:[ 0 5 9 13 0 ]
  //: joint g34 (P1) @(3, -87) /w:[ 12 14 -1 11 ]
  //: joint g28 (P0) @(73, -179) /w:[ 12 14 -1 11 ]
  //: joint g57 (P3) @(-103, 217) /w:[ 14 13 -1 16 ]
  //: output g46 (PG) @(432,151) /sn:0 /w:[ 1 ]
  and g11 (.I0(G0), .I1(P1), .Z(w8));   //: @(253,-86) /sn:0 /w:[ 7 13 0 ]
  //: input g5 (G2) @(-40,-205) /sn:0 /R:3 /w:[ 3 ]
  and g14 (.I0(G1), .I1(P2), .Z(w17));   //: @(260,42) /sn:0 /w:[ 7 5 0 ]
  and g61 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .I4(P3), .Z(w3));   //: @(236,111) /sn:0 /w:[ 13 0 0 0 0 0 ]
  or g19 (.I0(w2), .I1(G0), .Z(C1));   //: @(373,-170) /sn:0 /w:[ 1 3 0 ]
  or g21 (.I0(w11), .I1(w14), .I2(w17), .I3(G2), .Z(C3));   //: @(372,13) /sn:0 /w:[ 1 1 1 0 0 ]
  //: joint g32 (P1) @(3, -108) /w:[ 16 18 -1 15 ]
  or g20 (.I0(w5), .I1(w8), .I2(G1), .Z(C2));   //: @(368,-87) /sn:0 /w:[ 1 1 0 0 ]
  //: joint g63 (P2) @(-63, 114) /w:[ 1 2 -1 16 ]
  //: joint g38 (P1) @(3, -23) /w:[ 8 10 -1 7 ]
  and g15 (.I0(P0), .I1(P1), .I2(P2), .I3(P3), .Z(PG));   //: @(237,153) /sn:0 /w:[ 17 23 19 7 0 ]
  //: joint g43 (G1) @(27, 36) /w:[ 6 5 -1 8 ]
  //: input g0 (P0) @(73,-207) /sn:0 /R:3 /w:[ 15 ]
  //: joint g27 (C0) @(154, -182) /w:[ 8 10 -1 7 ]
  //: joint g48 (P1) @(3, 148) /w:[ 22 21 -1 24 ]
  //: joint g37 (P0) @(73, -28) /w:[ 4 6 -1 3 ]
  //: joint g62 (P3) @(-103, 120) /w:[ 1 2 -1 4 ]
  and g13 (.I0(G0), .I1(P1), .I2(P2), .Z(w14));   //: @(258,10) /sn:0 /w:[ 11 5 9 0 ]
  //: joint g53 (P2) @(-63, 184) /w:[ 22 21 -1 24 ]

endmodule

module CLA16_2(A, C4, PG, B, C0, GG, S);
//: interface  /sz:(140, 142) /bd:[ Ti0>A[15:0](37/140) Ti1>B[15:0](95/140) Li0>C0(61/142) Bo0<S[15:0](67/140) Ro0<C4(47/142) Ro1<PG(75/142) Ro2<GG(108/142) ]
input [15:0] B;    //: /sn:0 {0}(119,123)(352,123){1}
//: {2}(353,123)(574,123){3}
//: {4}(575,123)(798,123){5}
//: {6}(799,123)(1030,123){7}
//: {8}(1031,123)(1205,123){9}
input C0;    //: /sn:0 {0}(89,284)(149,284){1}
//: {2}(153,284)(176,284)(176,283)(274,283){3}
//: {4}(151,286)(151,429)(198,429){5}
output GG;    //: /sn:0 {0}(1082,490)(1082,460){1}
input [15:0] A;    //: /sn:0 {0}(120,88)(287,88){1}
//: {2}(288,88)(513,88){3}
//: {4}(514,88)(733,88){5}
//: {6}(734,88)(965,88){7}
//: {8}(966,88)(1203,88){9}
output PG;    //: /sn:0 {0}(1108,491)(1108,460){1}
output C4;    //: /sn:0 {0}(1190,431)(1160,431)(1160,432)(1150,432){1}
output [15:0] S;    //: /sn:0 /dp:1 {0}(1185,605)(1340,605){1}
wire [3:0] w6;    //: /sn:0 /dp:1 {0}(514,92)(514,224)(511,224)(511,234){1}
wire [3:0] w13;    //: /sn:0 {0}(569,234)(569,218)(575,218)(575,127){1}
wire [3:0] w7;    //: /sn:0 {0}(1179,590)(1018,590)(1018,330){1}
wire w25;    //: /sn:0 {0}(428,401)(428,284)(497,284){1}
wire [3:0] w3;    //: /sn:0 {0}(288,233)(288,92){1}
wire [3:0] w0;    //: /sn:0 {0}(1179,620)(358,620)(358,331){1}
wire w30;    //: /sn:0 {0}(768,401)(768,339)(757,339)(757,329){1}
wire w37;    //: /sn:0 {0}(731,329)(731,391)(737,391)(737,401){1}
wire w23;    //: /sn:0 {0}(270,401)(270,341)(299,341)(299,331){1}
wire w24;    //: /sn:0 {0}(299,401)(299,361)(324,361)(324,331){1}
wire w31;    //: /sn:0 {0}(852,401)(852,282)(934,282){1}
wire [3:0] w1;    //: /sn:0 {0}(353,127)(353,223)(346,223)(346,233){1}
wire w32;    //: /sn:0 {0}(955,401)(955,340)(959,340)(959,330){1}
wire w27;    //: /sn:0 {0}(535,401)(535,342)(547,342)(547,332){1}
wire w17;    //: /sn:0 {0}(522,332)(522,391)(508,391)(508,401){1}
wire w44;    //: /sn:0 {0}(984,330)(984,391)(987,391)(987,401){1}
wire w28;    //: /sn:0 {0}(643,401)(643,281)(705,281){1}
wire [3:0] w35;    //: /sn:0 {0}(780,231)(780,210)(799,210)(799,127){1}
wire [3:0] w11;    //: /sn:0 /dp:1 {0}(734,92)(734,210)(719,210)(719,231){1}
wire [3:0] w41;    //: /sn:0 {0}(1006,232)(1006,192)(1031,192)(1031,127){1}
wire [3:0] w2;    //: /sn:0 {0}(1179,610)(581,610)(581,332){1}
wire [3:0] w5;    //: /sn:0 {0}(1179,600)(793,600)(793,329){1}
wire [3:0] w40;    //: /sn:0 {0}(948,232)(948,192)(966,192)(966,92){1}
//: enddecls

  //: input g4 (A) @(118,88) /sn:0 /w:[ 0 ]
  tran g8(.Z(w6), .I(A[7:4]));   //: @(514,86) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  CLA_2 g3 (.B(w41), .A(w40), .C0(w31), .S(w7), .GG(w44), .PG(w32));   //: @(935, 233) /sz:(99, 96) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Bo1<0 Bo2<1 ]
  //: joint g16 (C0) @(151, 284) /w:[ 2 -1 1 4 ]
  //: output g17 (C4) @(1187,431) /sn:0 /w:[ 0 ]
  CLA_2 g2 (.B(w35), .A(w11), .C0(w28), .S(w5), .GG(w30), .PG(w37));   //: @(706, 232) /sz:(104, 96) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Bo0<1 Bo1<1 Bo2<0 ]
  CLA_2 g1 (.B(w13), .A(w6), .C0(w25), .S(w2), .GG(w27), .PG(w17));   //: @(498, 235) /sz:(99, 96) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Bo0<1 Bo1<1 Bo2<0 ]
  //: output g18 (PG) @(1108,488) /sn:0 /R:3 /w:[ 0 ]
  tran g10(.Z(w11), .I(A[11:8]));   //: @(734,86) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g6(.Z(w3), .I(A[3:0]));   //: @(288,86) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g7(.Z(w1), .I(B[3:0]));   //: @(353,121) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g9(.Z(w13), .I(B[7:4]));   //: @(575,121) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g12(.Z(w40), .I(A[15:12]));   //: @(966,86) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: input g5 (B) @(117,123) /sn:0 /w:[ 0 ]
  tran g11(.Z(w35), .I(B[11:8]));   //: @(799,121) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g14 (C0) @(87,284) /sn:0 /w:[ 0 ]
  //: output g19 (GG) @(1082,487) /sn:0 /R:3 /w:[ 0 ]
  concat g21 (.I0(w0), .I1(w2), .I2(w5), .I3(w7), .Z(S));   //: @(1184,605) /sn:0 /w:[ 0 0 0 0 0 ] /dr:0
  //: output g20 (S) @(1337,605) /sn:0 /w:[ 1 ]
  CLU_16 g15 (.G3(w44), .P3(w32), .G2(w30), .P2(w37), .G1(w27), .P1(w17), .G0(w24), .P0(w23), .C0(C0), .C3(w31), .C2(w28), .C1(w25), .GG(GG), .PG(PG), .C4(C4));   //: @(199, 402) /sz:(950, 57) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Ti3>1 Ti4>0 Ti5>1 Ti6>0 Ti7>0 Li0>5 To0<0 To1<0 To2<0 Bo0<1 Bo1<1 Ro0<1 ]
  CLA_2 g0 (.B(w1), .A(w3), .C0(C0), .S(w0), .GG(w24), .PG(w23));   //: @(275, 234) /sz:(99, 96) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>3 Bo0<1 Bo1<1 Bo2<1 ]
  tran g13(.Z(w41), .I(B[15:12]));   //: @(1031,121) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1

endmodule

module CLL(C1, P3, G3, P0, C3, C0, C4, P1, P2, G0, C2, G2, G1);
//: interface  /sz:(622, 40) /bd:[ Ti0>G0(67/622) Ti1>P0(100/622) Ti2>C1(152/622) Ti3>G1(232/622) Ti4>P1(261/622) Ti5>C2(323/622) Ti6>G2(384/622) Ti7>P2(412/622) Ti8>C3(477/622) Ti9>G3(554/622) Ti10>P3(584/622) Li0>C0(19/40) To0<C0(176/622) Ro0<C4(19/40) ]
input G2;    //: /sn:0 /dp:3 {0}(602,341)(140,341)(140,265)(120,265){1}
//: {2}(116,265)(51,265){3}
//: {4}(118,267)(118,461)(317,461){5}
input C0;    //: /sn:0 {0}(51,65)(205,65){1}
//: {2}(209,65)(401,65)(401,126)(403,126){3}
//: {4}(207,67)(207,155)(241,155){5}
//: {6}(245,155)(278,155)(278,179)(324,179){7}
//: {8}(243,157)(243,250)(249,250){9}
//: {10}(253,250)(326,250){11}
//: {12}(251,252)(251,353)(316,353){13}
input P1;    //: /sn:0 /dp:1 {0}(316,363)(242,363){1}
//: {2}(238,363)(221,363)(221,282){3}
//: {4}(223,280)(326,280){5}
//: {6}(219,280)(210,280)(210,262){7}
//: {8}(212,260)(326,260){9}
//: {10}(208,260)(201,260)(201,211){11}
//: {12}(203,209)(324,209){13}
//: {14}(199,209)(192,209)(192,182){15}
//: {16}(194,180)(264,180)(264,189)(324,189){17}
//: {18}(190,180)(52,180){19}
//: {20}(240,365)(240,399)(316,399){21}
output C3;    //: /sn:0 {0}(661,333)(623,333){1}
input G0;    //: /sn:0 {0}(52,140)(157,140){1}
//: {2}(161,140)(605,140){3}
//: {4}(159,142)(159,204)(168,204){5}
//: {6}(172,204)(324,204){7}
//: {8}(170,206)(170,275)(176,275){9}
//: {10}(180,275)(326,275){11}
//: {12}(178,277)(178,394)(316,394){13}
output C4;    //: /sn:0 /dp:1 {0}(621,423)(658,423){1}
output C2;    //: /sn:0 {0}(660,228)(623,228){1}
input P3;    //: /sn:0 {0}(316,436)(142,436)(142,411){1}
//: {2}(144,409)(316,409){3}
//: {4}(140,409)(109,409)(109,315){5}
//: {6}(111,313)(279,313)(279,373)(316,373){7}
//: {8}(107,313)(49,313){9}
input G1;    //: /sn:0 {0}(602,233)(104,233){1}
//: {2}(100,233)(71,233)(71,202)(51,202){3}
//: {4}(102,235)(102,299)(127,299){5}
//: {6}(131,299)(326,299){7}
//: {8}(129,301)(129,426)(316,426){9}
input G3;    //: /sn:0 /dp:1 {0}(317,466)(100,466)(100,333)(49,333){1}
input P0;    //: /sn:0 /dp:1 {0}(52,120)(176,120){1}
//: {2}(180,120)(371,120)(371,131)(403,131){3}
//: {4}(178,122)(178,184)(218,184){5}
//: {6}(222,184)(324,184){7}
//: {8}(220,186)(220,255)(227,255){9}
//: {10}(231,255)(326,255){11}
//: {12}(229,257)(229,358)(316,358){13}
output C1;    //: /sn:0 {0}(664,138)(626,138){1}
input P2;    //: /sn:0 {0}(316,404)(233,404){1}
//: {2}(229,404)(210,404)(210,370){3}
//: {4}(212,368)(316,368){5}
//: {6}(208,368)(201,368)(201,306){7}
//: {8}(203,304)(326,304){9}
//: {10}(199,304)(185,304)(185,287){11}
//: {12}(187,285)(326,285){13}
//: {14}(183,285)(154,285)(154,245){15}
//: {16}(156,243)(288,243)(288,265)(326,265){17}
//: {18}(152,243)(52,243){19}
//: {20}(231,406)(231,431)(316,431){21}
wire w7;    //: /sn:0 /dp:1 {0}(602,331)(582,331)(582,280)(347,280){1}
wire w4;    //: /sn:0 /dp:1 {0}(602,228)(559,228)(559,207)(345,207){1}
wire w42;    //: /sn:0 {0}(602,336)(574,336)(574,302)(347,302){1}
wire w24;    //: /sn:0 {0}(337,363)(590,363)(590,416)(600,416){1}
wire w8;    //: /sn:0 {0}(424,129)(595,129)(595,135)(605,135){1}
wire w27;    //: /sn:0 {0}(337,401)(584,401)(584,421)(600,421){1}
wire w33;    //: /sn:0 {0}(338,464)(590,464)(590,431)(600,431){1}
wire w41;    //: /sn:0 {0}(600,426)(572,426)(572,431)(337,431){1}
wire w2;    //: /sn:0 {0}(345,184)(592,184)(592,223)(602,223){1}
wire w15;    //: /sn:0 {0}(347,257)(592,257)(592,326)(602,326){1}
//: enddecls

  //: joint g44 (G0) @(178, 275) /w:[ 10 -1 9 12 ]
  and g8 (.I0(C0), .I1(P0), .Z(w8));   //: @(414,129) /sn:0 /w:[ 3 3 0 ]
  //: output g4 (C1) @(661,138) /sn:0 /w:[ 0 ]
  //: joint g47 (P3) @(109, 313) /w:[ 6 -1 8 5 ]
  //: input g16 (P3) @(47,313) /sn:0 /w:[ 9 ]
  or g3 (.I0(w24), .I1(w27), .I2(w41), .I3(w33), .Z(C4));   //: @(611,423) /sn:0 /w:[ 1 1 0 1 0 ]
  and g26 (.I0(G2), .I1(G3), .Z(w33));   //: @(328,464) /sn:0 /w:[ 5 0 0 ]
  //: input g17 (G3) @(47,333) /sn:0 /w:[ 1 ]
  or g2 (.I0(w15), .I1(w7), .I2(w42), .I3(G2), .Z(C3));   //: @(613,333) /sn:0 /w:[ 1 0 0 0 1 ]
  //: joint g30 (G0) @(159, 140) /w:[ 2 -1 1 4 ]
  and g23 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .I4(P3), .Z(w24));   //: @(327,363) /sn:0 /w:[ 13 13 0 5 7 0 ]
  //: joint g39 (P2) @(185, 285) /w:[ 12 -1 14 11 ]
  and g24 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w27));   //: @(327,401) /sn:0 /w:[ 13 21 0 3 0 ]
  or g1 (.I0(w2), .I1(w4), .I2(G1), .Z(C2));   //: @(613,228) /sn:0 /w:[ 1 0 0 1 ]
  //: joint g29 (P0) @(178, 120) /w:[ 2 -1 1 4 ]
  and g18 (.I0(C0), .I1(P0), .I2(P1), .Z(w2));   //: @(335,184) /sn:0 /w:[ 7 7 17 0 ]
  and g25 (.I0(G1), .I1(P2), .I2(P3), .Z(w41));   //: @(327,431) /sn:0 /w:[ 9 21 0 1 ]
  //: input g10 (P0) @(50,120) /sn:0 /w:[ 0 ]
  //: joint g49 (P2) @(231, 404) /w:[ 1 -1 2 20 ]
  //: joint g50 (P3) @(142, 409) /w:[ 2 -1 4 1 ]
  //: output g6 (C3) @(658,333) /sn:0 /w:[ 0 ]
  //: joint g35 (G0) @(170, 204) /w:[ 6 -1 5 8 ]
  //: input g9 (C0) @(49,65) /sn:0 /w:[ 0 ]
  //: output g7 (C4) @(655,423) /sn:0 /w:[ 1 ]
  //: joint g31 (P1) @(192, 180) /w:[ 16 -1 18 15 ]
  and g22 (.I0(G1), .I1(P2), .Z(w42));   //: @(337,302) /sn:0 /w:[ 7 9 1 ]
  //: joint g45 (P1) @(240, 363) /w:[ 1 -1 2 20 ]
  //: joint g41 (P0) @(229, 255) /w:[ 10 -1 9 12 ]
  //: joint g36 (P1) @(210, 260) /w:[ 8 -1 10 7 ]
  //: joint g33 (P0) @(220, 184) /w:[ 6 -1 5 8 ]
  //: joint g42 (P1) @(221, 280) /w:[ 4 -1 6 3 ]
  //: joint g40 (C0) @(251, 250) /w:[ 10 -1 9 12 ]
  //: input g12 (P1) @(50,180) /sn:0 /w:[ 19 ]
  //: joint g46 (P2) @(210, 368) /w:[ 4 -1 6 3 ]
  //: joint g34 (P1) @(201, 209) /w:[ 12 -1 14 11 ]
  //: joint g28 (C0) @(207, 65) /w:[ 2 -1 1 4 ]
  //: input g14 (P2) @(50,243) /sn:0 /w:[ 19 ]
  //: input g11 (G0) @(50,140) /sn:0 /w:[ 0 ]
  //: output g5 (C2) @(657,228) /sn:0 /w:[ 0 ]
  and g21 (.I0(G0), .I1(P1), .I2(P2), .Z(w7));   //: @(337,280) /sn:0 /w:[ 11 5 13 1 ]
  and g19 (.I0(G0), .I1(P1), .Z(w4));   //: @(335,207) /sn:0 /w:[ 7 13 1 ]
  //: joint g32 (C0) @(243, 155) /w:[ 6 -1 5 8 ]
  and g20 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .Z(w15));   //: @(337,257) /sn:0 /w:[ 11 11 9 17 0 ]
  //: joint g43 (P2) @(201, 304) /w:[ 8 -1 10 7 ]
  //: joint g38 (G1) @(102, 233) /w:[ 1 -1 2 4 ]
  //: input g15 (G2) @(49,265) /sn:0 /w:[ 3 ]
  or g0 (.I0(w8), .I1(G0), .Z(C1));   //: @(616,138) /sn:0 /w:[ 1 3 1 ]
  //: joint g48 (G1) @(129, 299) /w:[ 6 -1 5 8 ]
  //: joint g27 (G2) @(118, 265) /w:[ 1 -1 2 4 ]
  //: joint g37 (P2) @(154, 243) /w:[ 16 -1 18 15 ]
  //: input g13 (G1) @(49,202) /sn:0 /w:[ 3 ]

endmodule

module CLL_2(C0, P2, P1, GG, G1, C1, C2, G0, C3, P3, G3, PG, G2, P0);
//: interface  /sz:(40, 40) /bd:[ ]
input G2;    //: /sn:0 {0}(367,-6)(309,-6)(309,36)(-99,36){1}
//: {2}(-101,34)(-101,-231){3}
//: {4}(-101,38)(-101,213)(74,213)(74,222)(247,222){5}
input C0;    //: /sn:0 /dp:7 {0}(235,-145)(137,-145)(137,-151)(85,-151){1}
//: {2}(83,-153)(83,-203){3}
//: {4}(85,-205)(142,-205)(142,-217)(236,-217){5}
//: {6}(83,-207)(83,-237){7}
//: {8}(83,-149)(83,-65)(138,-65)(138,-57)(243,-57){9}
output GG;    //: /sn:0 {0}(392,178)(412,178){1}
input P1;    //: /sn:0 {0}(244,125)(-5,125)(-5,117)(-56,117){1}
//: {2}(-58,115)(-58,-20){3}
//: {4}(-56,-22)(95,-22)(95,-18)(241,-18){5}
//: {6}(-58,-24)(-58,-52){7}
//: {8}(-56,-54)(-3,-54)(-3,-47)(243,-47){9}
//: {10}(-58,-56)(-58,-101){11}
//: {12}(-56,-103)(62,-103)(62,-112)(236,-112){13}
//: {14}(-58,-105)(-58,-137){15}
//: {16}(-56,-139)(92,-139)(92,-135)(235,-135){17}
//: {18}(-58,-141)(-58,-232){19}
//: {20}(-58,119)(-58,149)(146,149)(146,157)(246,157){21}
output C3;    //: /sn:0 {0}(388,-14)(402,-14)(402,-7)(412,-7){1}
output PG;    //: /sn:0 {0}(265,127)(401,127)(401,128)(411,128){1}
input G0;    //: /sn:0 {0}(39,-234)(39,-197){1}
//: {2}(41,-195)(121,-195)(121,-197)(346,-197){3}
//: {4}(39,-193)(39,-122){5}
//: {6}(41,-120)(150,-120)(150,-117)(236,-117){7}
//: {8}(39,-118)(39,-28){9}
//: {10}(41,-26)(153,-26)(153,-23)(241,-23){11}
//: {12}(39,-24)(39,152)(246,152){13}
output C2;    //: /sn:0 {0}(378,-110)(402,-110)(402,-108)(412,-108){1}
input P3;    //: /sn:0 {0}(247,197)(-114,197)(-114,190)(-165,190){1}
//: {2}(-167,188)(-167,161){3}
//: {4}(-165,159)(-115,159)(-115,167)(246,167){5}
//: {6}(-167,157)(-167,134){7}
//: {8}(-165,132)(24,132)(24,135)(244,135){9}
//: {10}(-167,130)(-167,-230){11}
//: {12}(-167,192)(-167,219)(32,219)(32,227)(247,227){13}
input G1;    //: /sn:0 {0}(357,-105)(183,-105)(183,-112)(-32,-112){1}
//: {2}(-34,-114)(-34,-234){3}
//: {4}(-34,-110)(-34,3){5}
//: {6}(-32,5)(20,5)(20,11)(243,11){7}
//: {8}(-34,7)(-34,187)(247,187){9}
input G3;    //: /sn:0 /dp:1 {0}(-183,-229)(-183,252)(303,252)(303,198)(331,198)(331,186)(371,186){1}
input P0;    //: /sn:0 /dp:11 {0}(243,-52)(141,-52)(141,-56)(14,-56){1}
//: {2}(12,-58)(12,-140){3}
//: {4}(14,-142)(66,-142)(66,-140)(235,-140){5}
//: {6}(12,-144)(12,-205){7}
//: {8}(14,-207)(138,-207)(138,-212)(236,-212){9}
//: {10}(12,-209)(12,-233){11}
//: {12}(12,-54)(12,113)(138,113)(138,120)(244,120){13}
output C1;    //: /sn:0 {0}(367,-199)(402,-199)(402,-191)(412,-191){1}
input P2;    //: /sn:0 {0}(246,162)(-72,162)(-72,156)(-122,156){1}
//: {2}(-124,154)(-124,129){3}
//: {4}(-122,127)(-46,127)(-46,99)(65,99)(65,130)(244,130){5}
//: {6}(-124,125)(-124,16){7}
//: {8}(-122,14)(-70,14)(-70,16)(243,16){9}
//: {10}(-124,12)(-124,-16){11}
//: {12}(-122,-18)(-70,-18)(-70,-13)(241,-13){13}
//: {14}(-124,-20)(-124,-43){15}
//: {16}(-122,-45)(54,-45)(54,-42)(243,-42){17}
//: {18}(-124,-47)(-124,-230){19}
//: {20}(-124,158)(-124,184)(146,184)(146,192)(247,192){21}
wire w29;    //: /sn:0 {0}(268,225)(352,225)(352,196)(361,196)(361,181)(371,181){1}
wire w23;    //: /sn:0 {0}(267,159)(361,159)(361,176)(371,176){1}
wire w8;    //: /sn:0 {0}(257,-114)(347,-114)(347,-110)(357,-110){1}
wire w17;    //: /sn:0 {0}(264,14)(357,14)(357,-11)(367,-11){1}
wire w14;    //: /sn:0 {0}(262,-18)(357,-18)(357,-16)(367,-16){1}
wire w2;    //: /sn:0 {0}(257,-214)(345,-214)(345,-202)(346,-202){1}
wire w11;    //: /sn:0 {0}(264,-50)(356,-50)(356,-21)(367,-21){1}
wire w5;    //: /sn:0 {0}(256,-140)(295,-140)(295,-125)(340,-125)(340,-115)(357,-115){1}
wire w26;    //: /sn:0 {0}(268,192)(304,192)(304,171)(371,171){1}
//: enddecls

  //: joint g44 (P2) @(-124, 14) /w:[ 8 10 -1 7 ]
  //: input g8 (C0) @(83,-239) /sn:0 /R:3 /w:[ 7 ]
  //: input g4 (P2) @(-124,-232) /sn:0 /R:3 /w:[ 19 ]
  and g16 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w23));   //: @(257,159) /sn:0 /w:[ 13 21 0 5 0 ]
  //: input g3 (P1) @(-58,-234) /sn:0 /R:3 /w:[ 19 ]
  //: output g26 (GG) @(409,178) /sn:0 /w:[ 1 ]
  and g17 (.I0(G1), .I1(P2), .I2(P3), .Z(w26));   //: @(258,192) /sn:0 /w:[ 9 21 0 0 ]
  //: input g2 (G1) @(-34,-236) /sn:0 /R:3 /w:[ 3 ]
  //: joint g30 (C0) @(83, -151) /w:[ 1 2 -1 8 ]
  //: output g23 (C1) @(409,-191) /sn:0 /w:[ 1 ]
  //: output g24 (C2) @(409,-108) /sn:0 /w:[ 1 ]
  //: joint g39 (P2) @(-124, -45) /w:[ 16 18 -1 15 ]
  //: input g1 (G0) @(39,-236) /sn:0 /R:3 /w:[ 0 ]
  //: joint g29 (G0) @(39, -195) /w:[ 2 1 -1 4 ]
  and g18 (.I0(G2), .I1(P3), .Z(w29));   //: @(258,225) /sn:0 /w:[ 5 13 0 ]
  //: output g25 (C3) @(409,-7) /sn:0 /w:[ 1 ]
  and g10 (.I0(C0), .I1(P0), .I2(P1), .Z(w5));   //: @(246,-140) /sn:0 /w:[ 0 5 17 0 ]
  //: joint g49 (P2) @(-124, 127) /w:[ 4 6 -1 3 ]
  //: input g6 (P3) @(-167,-232) /sn:0 /R:3 /w:[ 11 ]
  //: joint g50 (P3) @(-167, 132) /w:[ 8 10 -1 7 ]
  //: joint g35 (G1) @(-34, -112) /w:[ 1 2 -1 4 ]
  and g9 (.I0(C0), .I1(P0), .Z(w2));   //: @(247,-214) /sn:0 /w:[ 5 9 0 ]
  //: input g7 (G3) @(-183,-231) /sn:0 /R:3 /w:[ 0 ]
  or g22 (.I0(w26), .I1(w23), .I2(w29), .I3(G3), .Z(GG));   //: @(382,178) /sn:0 /w:[ 1 1 1 1 0 ]
  //: joint g31 (P0) @(12, -142) /w:[ 4 6 -1 3 ]
  //: joint g33 (G0) @(39, -120) /w:[ 6 5 -1 8 ]
  //: joint g45 (G2) @(-101, 36) /w:[ 1 2 -1 4 ]
  //: joint g54 (P3) @(-167, 159) /w:[ 4 6 -1 3 ]
  //: joint g41 (P1) @(-58, -22) /w:[ 4 6 -1 3 ]
  //: joint g40 (G0) @(39, -26) /w:[ 10 9 -1 12 ]
  //: joint g42 (P2) @(-124, -18) /w:[ 12 14 -1 11 ]
  and g12 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .Z(w11));   //: @(254,-50) /sn:0 /w:[ 9 0 9 17 0 ]
  //: output g46 (PG) @(408,128) /sn:0 /w:[ 1 ]
  //: joint g57 (P3) @(-167, 190) /w:[ 1 2 -1 12 ]
  //: joint g28 (P0) @(12, -207) /w:[ 8 10 -1 7 ]
  //: joint g34 (P1) @(-58, -103) /w:[ 12 14 -1 11 ]
  and g14 (.I0(G1), .I1(P2), .Z(w17));   //: @(254,14) /sn:0 /w:[ 7 9 0 ]
  //: input g5 (G2) @(-101,-233) /sn:0 /R:3 /w:[ 3 ]
  and g11 (.I0(G0), .I1(P1), .Z(w8));   //: @(247,-114) /sn:0 /w:[ 7 13 0 ]
  or g21 (.I0(w11), .I1(w14), .I2(w17), .I3(G2), .Z(C3));   //: @(378,-14) /sn:0 /w:[ 1 1 1 0 0 ]
  or g19 (.I0(w2), .I1(G0), .Z(C1));   //: @(357,-199) /sn:0 /w:[ 1 3 0 ]
  or g20 (.I0(w5), .I1(w8), .I2(G1), .Z(C2));   //: @(368,-110) /sn:0 /w:[ 1 1 0 0 ]
  //: joint g32 (P1) @(-58, -139) /w:[ 16 18 -1 15 ]
  //: input g0 (P0) @(12,-235) /sn:0 /R:3 /w:[ 11 ]
  //: joint g43 (G1) @(-34, 5) /w:[ 6 5 -1 8 ]
  and g15 (.I0(P0), .I1(P1), .I2(P2), .I3(P3), .Z(PG));   //: @(255,127) /sn:0 /w:[ 13 0 5 9 0 ]
  //: joint g38 (P1) @(-58, -54) /w:[ 8 10 -1 7 ]
  //: joint g48 (P1) @(-58, 117) /w:[ 1 2 -1 20 ]
  //: joint g27 (C0) @(83, -205) /w:[ 4 6 -1 3 ]
  //: joint g37 (P0) @(12, -56) /w:[ 1 2 -1 12 ]
  //: joint g53 (P2) @(-124, 156) /w:[ 1 2 -1 20 ]
  and g13 (.I0(G0), .I1(P1), .I2(P2), .Z(w14));   //: @(252,-18) /sn:0 /w:[ 11 5 13 0 ]

endmodule

module PFA(A, Pi, Ci, S, Gi, B);
//: interface  /sz:(100, 97) /bd:[ Ti0>B(50/100) Ti1>A(14/100) Li0>Ci(46/97) Bo0<Gi(61/100) Ro0<Pi(67/97) Ro1<S(32/97) ]
input B;    //: /sn:0 {0}(184,223)(195,223){1}
//: {2}(199,223)(226,223)(226,207)(234,207){3}
//: {4}(197,225)(197,256){5}
//: {6}(199,258)(308,258){7}
//: {8}(197,260)(197,293)(309,293){9}
output Gi;    //: /sn:0 /dp:1 {0}(330,291)(354,291){1}
input A;    //: /sn:0 {0}(186,202)(214,202){1}
//: {2}(218,202)(234,202){3}
//: {4}(216,204)(216,251){5}
//: {6}(218,253)(308,253){7}
//: {8}(216,255)(216,288)(309,288){9}
output Pi;    //: /sn:0 /dp:1 {0}(329,256)(351,256){1}
input Ci;    //: /sn:0 /dp:1 {0}(305,227)(274,227)(274,241)(187,241){1}
output S;    //: /sn:0 {0}(358,225)(326,225){1}
wire w11;    //: /sn:0 {0}(255,205)(295,205)(295,222)(305,222){1}
//: enddecls

  //: input g4 (A) @(184,202) /sn:0 /w:[ 0 ]
  //: output g8 (Pi) @(348,256) /sn:0 /w:[ 1 ]
  xor g3 (.I0(A), .I1(B), .Z(w11));   //: @(245,205) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  xor g2 (.I0(w11), .I1(Ci), .Z(S));   //: @(316,225) /sn:0 /delay:" 2" /w:[ 1 0 1 ]
  or g1 (.I0(A), .I1(B), .Z(Pi));   //: @(319,256) /sn:0 /w:[ 7 7 0 ]
  //: joint g10 (A) @(216, 202) /w:[ 2 -1 1 4 ]
  //: input g6 (Ci) @(185,241) /sn:0 /w:[ 1 ]
  //: output g7 (S) @(355,225) /sn:0 /w:[ 0 ]
  //: output g9 (Gi) @(351,291) /sn:0 /w:[ 1 ]
  //: joint g12 (A) @(216, 253) /w:[ 6 5 -1 8 ]
  //: input g5 (B) @(182,223) /sn:0 /w:[ 0 ]
  //: joint g11 (B) @(197, 223) /w:[ 2 -1 1 4 ]
  and g0 (.I0(A), .I1(B), .Z(Gi));   //: @(320,291) /sn:0 /w:[ 9 9 0 ]
  //: joint g13 (B) @(197, 258) /w:[ 6 5 -1 8 ]

endmodule

module main;    //: root_module
wire w88;    //: /sn:0 {0}(-148,31)(-246,31)(-246,89)(-274,89){1}
wire [3:0] w72;    //: /sn:0 /dp:1 {0}(184,260)(184,318)(30,318){1}
wire w62;    //: /sn:0 {0}(-134,137)(-110,137){1}
wire w109;    //: /sn:0 {0}(95,34)(143,34)(143,102)(221,102){1}
wire w101;    //: /sn:0 {0}(95,-46)(183,-46)(183,-122)(220,-122){1}
wire w82;    //: /sn:0 /dp:1 {0}(-148,81)(-196,81)(-196,230)(-274,230){1}
wire [3:0] w71;    //: /sn:0 {0}(129,259)(129,298)(30,298){1}
wire w112;    //: /sn:0 {0}(95,64)(118,64)(118,187)(221,187){1}
wire w66;    //: /sn:0 {0}(69,123)(32,123){1}
wire [15:0] w12;    //: /sn:0 /dp:1 {0}(-72,75)(-72,6)(-142,6){1}
wire [15:0] w63;    //: /sn:0 /dp:1 {0}(24,303)(-42,303)(-42,219){1}
wire [3:0] w70;    //: /sn:0 {0}(100,259)(100,288)(30,288){1}
wire w111;    //: /sn:0 {0}(95,54)(125,54)(125,158)(221,158){1}
wire w91;    //: /sn:0 {0}(-148,1)(-266,1)(-266,6)(-275,6){1}
wire w108;    //: /sn:0 {0}(95,24)(152,24)(152,74)(221,74){1}
wire w86;    //: /sn:0 {0}(95,-86)(142,-86)(142,-235)(220,-235){1}
wire w106;    //: /sn:0 {0}(95,4)(172,4)(172,17)(221,17){1}
wire w104;    //: /sn:0 {0}(95,-16)(211,-16)(211,-37)(220,-37){1}
wire w68;    //: /sn:0 {0}(56,182)(41,182)(41,184)(32,184){1}
wire w110;    //: /sn:0 {0}(95,44)(135,44)(135,130)(221,130){1}
wire w103;    //: /sn:0 {0}(95,-26)(203,-26)(203,-66)(220,-66){1}
wire w98;    //: /sn:0 {0}(-148,-69)(-172,-69)(-172,-192)(-275,-192){1}
wire w95;    //: /sn:0 {0}(-148,-39)(-197,-39)(-197,-107)(-275,-107){1}
wire w89;    //: /sn:0 {0}(-148,21)(-257,21)(-257,61)(-274,61){1}
wire [15:0] w113;    //: /sn:0 /dp:1 {0}(89,-11)(-14,-11)(-14,75){1}
wire w80;    //: /sn:0 {0}(220,-150)(175,-150)(175,-56)(95,-56){1}
wire w67;    //: /sn:0 {0}(59,150)(42,150)(42,151)(32,151){1}
wire [3:0] w69;    //: /sn:0 /dp:1 {0}(156,259)(156,308)(30,308){1}
wire w105;    //: /sn:0 {0}(95,-6)(212,-6)(212,-11)(221,-11){1}
wire w90;    //: /sn:0 {0}(-148,11)(-265,11)(-265,32)(-274,32){1}
wire w85;    //: /sn:0 {0}(-148,61)(-215,61)(-215,174)(-274,174){1}
wire w83;    //: /sn:0 /dp:1 {0}(-148,71)(-209,71)(-209,202)(-274,202){1}
wire w102;    //: /sn:0 {0}(95,-36)(192,-36)(192,-94)(220,-94){1}
wire w94;    //: /sn:0 {0}(-148,-29)(-206,-29)(-206,-79)(-275,-79){1}
wire w92;    //: /sn:0 {0}(-148,-9)(-226,-9)(-226,-22)(-275,-22){1}
wire w87;    //: /sn:0 {0}(-148,41)(-237,41)(-237,117)(-274,117){1}
wire w107;    //: /sn:0 {0}(95,14)(161,14)(161,45)(221,45){1}
wire w100;    //: /sn:0 {0}(95,-66)(161,-66)(161,-179)(220,-179){1}
wire w99;    //: /sn:0 {0}(95,-76)(155,-76)(155,-207)(220,-207){1}
wire w97;    //: /sn:0 {0}(-148,-59)(-179,-59)(-179,-163)(-275,-163){1}
wire w96;    //: /sn:0 {0}(-148,-49)(-189,-49)(-189,-135)(-275,-135){1}
wire w93;    //: /sn:0 {0}(-148,-19)(-215,-19)(-215,-50)(-275,-50){1}
wire w79;    //: /sn:0 {0}(-274,145)(-229,145)(-229,51)(-148,51){1}
//: enddecls

  concat g75 (.I0(w82), .I1(w83), .I2(w85), .I3(w79), .I4(w87), .I5(w88), .I6(w89), .I7(w90), .I8(w91), .I9(w92), .I10(w93), .I11(w94), .I12(w95), .I13(w96), .I14(w97), .I15(w98), .Z(w12));   //: @(-143,6) /sn:0 /w:[ 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0
  //: switch g90 (w110) @(239,130) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: switch g92 (w109) @(239,102) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: switch g91 (w107) @(239,45) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: switch g74 (w82) @(-291,230) /sn:0 /w:[ 1 ] /st:1
  //: switch g86 (w100) @(238,-179) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: switch g77 (w86) @(238,-235) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: switch g60 (w97) @(-292,-163) /sn:0 /w:[ 1 ] /st:1
  //: switch g82 (w80) @(238,-150) /sn:0 /R:2 /w:[ 0 ] /st:1
  //: switch g70 (w87) @(-291,117) /sn:0 /w:[ 1 ] /st:1
  led g94 (.I(w69));   //: @(156,252) /sn:0 /w:[ 0 ] /type:1
  //: switch g65 (w92) @(-292,-22) /sn:0 /w:[ 1 ] /st:1
  //: switch g64 (w94) @(-292,-79) /sn:0 /w:[ 1 ] /st:1
  //: switch g72 (w79) @(-291,145) /sn:0 /w:[ 0 ] /st:1
  //: switch g73 (w83) @(-291,202) /sn:0 /w:[ 1 ] /st:1
  //: switch g68 (w90) @(-291,32) /sn:0 /w:[ 1 ] /st:1
  //: switch g58 (w62) @(-151,137) /sn:0 /w:[ 0 ] /st:1
  led g56 (.I(w67));   //: @(66,150) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: switch g71 (w85) @(-291,174) /sn:0 /w:[ 1 ] /st:1
  //: switch g59 (w98) @(-292,-192) /sn:0 /w:[ 1 ] /st:1
  //: switch g87 (w103) @(238,-66) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: switch g85 (w112) @(239,187) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: switch g67 (w89) @(-291,61) /sn:0 /w:[ 1 ] /st:1
  //: switch g83 (w104) @(238,-37) /sn:0 /R:2 /w:[ 1 ] /st:1
  CLA16_2 g54 (.B(w113), .A(w12), .C0(w62), .S(w63), .GG(w68), .PG(w67), .C4(w66));   //: @(-109, 76) /sz:(140, 142) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Bo0<1 Ro0<1 Ro1<1 Ro2<1 ]
  //: switch g81 (w108) @(239,74) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: switch g69 (w88) @(-291,89) /sn:0 /w:[ 1 ] /st:1
  //: switch g66 (w91) @(-292,6) /sn:0 /w:[ 1 ] /st:1
  led g57 (.I(w68));   //: @(63,182) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: switch g84 (w99) @(238,-207) /sn:0 /R:2 /w:[ 1 ] /st:1
  led g96 (.I(w71));   //: @(129,252) /sn:0 /w:[ 0 ] /type:1
  //: switch g61 (w96) @(-292,-135) /sn:0 /w:[ 1 ] /st:1
  //: switch g79 (w101) @(238,-122) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: switch g78 (w111) @(239,158) /sn:0 /R:2 /w:[ 1 ] /st:1
  led g97 (.I(w72));   //: @(184,253) /sn:0 /w:[ 0 ] /type:1
  concat g93 (.I0(w70), .I1(w71), .I2(w69), .I3(w72), .Z(w63));   //: @(25,303) /sn:0 /R:2 /w:[ 1 1 1 1 0 ] /dr:0
  //: switch g63 (w93) @(-292,-50) /sn:0 /w:[ 1 ] /st:1
  //: switch g89 (w105) @(239,-11) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: switch g62 (w95) @(-292,-107) /sn:0 /w:[ 1 ] /st:1
  led g95 (.I(w70));   //: @(100,252) /sn:0 /w:[ 0 ] /type:1
  //: switch g88 (w102) @(238,-94) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: switch g80 (w106) @(239,17) /sn:0 /R:2 /w:[ 1 ] /st:1
  led g55 (.I(w66));   //: @(76,123) /sn:0 /R:3 /w:[ 0 ] /type:0
  concat g76 (.I0(w86), .I1(w99), .I2(w100), .I3(w80), .I4(w101), .I5(w102), .I6(w103), .I7(w104), .I8(w105), .I9(w106), .I10(w107), .I11(w108), .I12(w109), .I13(w110), .I14(w111), .I15(w112), .Z(w113));   //: @(90,-11) /sn:0 /R:2 /w:[ 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /dr:0

endmodule

module CLA(A, C4, B, S, C0);
//: interface  /sz:(122, 98) /bd:[ Ti0>A[3:0](23/122) Ti1>B[3:0](88/122) Li0>C0(46/98) Bo0<S[3:0](66/122) Ro0<C4(52/98) ]
input [3:0] B;    //: /sn:0 /dp:1 {0}(40,86)(137,86){1}
//: {2}(138,86)(301,86){3}
//: {4}(302,86)(459,86){5}
//: {6}(460,86)(621,86){7}
//: {8}(622,86)(726,86){9}
input C0;    //: /sn:0 {0}(30,251)(40,251){1}
//: {2}(44,251)(52,251)(52,215)(87,215){3}
//: {4}(42,253)(42,372)(61,372){5}
input [3:0] A;    //: /sn:0 {0}(42,61)(101,61){1}
//: {2}(102,61)(138,61)(138,61)(265,61){3}
//: {4}(266,61)(423,61){5}
//: {6}(424,61)(585,61){7}
//: {8}(586,61)(732,61){9}
output C4;    //: /sn:0 {0}(739,372)(685,372){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(760,529)(739,529){1}
wire w13;    //: /sn:0 {0}(424,170)(424,65){1}
wire w6;    //: /sn:0 {0}(302,170)(302,90){1}
wire w7;    //: /sn:0 {0}(266,170)(266,65){1}
wire w34;    //: /sn:0 /dp:1 {0}(549,352)(549,220)(571,220){1}
wire w3;    //: /sn:0 /dp:1 {0}(733,534)(381,534)(381,203)(353,203){1}
wire w0;    //: /sn:0 {0}(138,168)(138,90){1}
wire w29;    //: /sn:0 /dp:1 {0}(321,352)(321,294)(368,294)(368,238)(353,238){1}
wire w19;    //: /sn:0 {0}(586,173)(586,65){1}
wire w18;    //: /sn:0 {0}(622,173)(622,90){1}
wire w12;    //: /sn:0 {0}(460,170)(460,90){1}
wire w10;    //: /sn:0 {0}(733,514)(705,514)(705,206)(673,206){1}
wire w21;    //: /sn:0 {0}(595,272)(595,352){1}
wire w31;    //: /sn:0 /dp:1 {0}(385,352)(385,217)(409,217){1}
wire w1;    //: /sn:0 {0}(102,168)(102,65){1}
wire w32;    //: /sn:0 /dp:1 {0}(471,352)(471,296)(525,296)(525,244)(511,244){1}
wire w8;    //: /sn:0 {0}(733,524)(541,524)(541,218)(511,218){1}
wire w27;    //: /sn:0 /dp:1 {0}(112,352)(112,267){1}
wire w28;    //: /sn:0 {0}(229,352)(229,217)(251,217){1}
wire w35;    //: /sn:0 /dp:1 {0}(638,352)(638,301)(688,301)(688,241)(673,241){1}
wire w2;    //: /sn:0 {0}(733,544)(212,544)(212,201)(189,201){1}
wire w15;    //: /sn:0 {0}(433,269)(433,352){1}
wire w26;    //: /sn:0 /dp:1 {0}(137,352)(137,320)(201,320)(201,236)(189,236){1}
wire w9;    //: /sn:0 {0}(278,269)(278,352){1}
//: enddecls

  tran g8(.Z(w7), .I(A[1]));   //: @(266,59) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: input g4 (A) @(40,61) /sn:0 /w:[ 0 ]
  //: joint g16 (C0) @(42, 251) /w:[ 2 -1 1 4 ]
  PFA g3 (.A(w19), .B(w18), .Ci(w34), .Gi(w21), .S(w10), .Pi(w35));   //: @(572, 174) /sz:(100, 97) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<1 Ro1<1 ]
  //: output g17 (C4) @(736,372) /sn:0 /w:[ 0 ]
  PFA g2 (.A(w13), .B(w12), .Ci(w31), .Gi(w15), .S(w8), .Pi(w32));   //: @(410, 171) /sz:(100, 97) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<1 Ro1<1 ]
  PFA g1 (.A(w7), .B(w6), .Ci(w28), .Gi(w9), .S(w3), .Pi(w29));   //: @(252, 171) /sz:(100, 97) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<1 Ro1<1 ]
  concat g18 (.I0(w2), .I1(w3), .I2(w8), .I3(w10), .Z(S));   //: @(738,529) /sn:0 /w:[ 0 0 0 0 1 ] /dr:0
  tran g10(.Z(w13), .I(A[2]));   //: @(424,59) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g6(.Z(w1), .I(A[0]));   //: @(102,59) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g7(.Z(w0), .I(B[0]));   //: @(138,84) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g9(.Z(w6), .I(B[1]));   //: @(302,84) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g12(.Z(w19), .I(A[3]));   //: @(586,59) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  CLL g14 (.P3(w21), .G3(w35), .P2(w15), .G2(w32), .P1(w9), .G1(w29), .P0(w27), .G0(w26), .C0(C0), .C3(w34), .C2(w31), .C1(w28), .C4(C4));   //: @(62, 353) /sz:(622, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>1 Ti3>0 Ti4>1 Ti5>0 Ti6>0 Ti7>0 Li0>5 To0<0 To1<0 To2<0 Ro0<1 ]
  tran g11(.Z(w12), .I(B[2]));   //: @(460,84) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g5 (B) @(38,86) /sn:0 /w:[ 0 ]
  //: output g19 (S) @(757,529) /sn:0 /w:[ 0 ]
  //: input g15 (C0) @(28,251) /sn:0 /w:[ 0 ]
  PFA g0 (.A(w1), .B(w0), .Ci(C0), .Gi(w27), .S(w2), .Pi(w26));   //: @(88, 169) /sz:(100, 97) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>3 Bo0<1 Ro0<1 Ro1<1 ]
  tran g13(.Z(w18), .I(B[3]));   //: @(622,84) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1

endmodule
