//: version "1.8.7"

module main;    //: root_module
input A0;    //: /sn:0 {0}(242,211)(258,211)(258,213)(279,213){1}
output C0;    //: /sn:0 {0}(515,277)(477,277)(477,278)(464,278){1}
output S0;    //: /sn:0 {0}(513,224)(464,224){1}
input B0;    //: /sn:0 {0}(246,275)(277,275)(277,276)(279,276){1}
//: enddecls

  HalfAdder g8 (.B(B0), .A(A0), .C(C0), .S(S0));   //: @(280, 185) /sz:(183, 127) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<1 ]
  //: input g10 (B0) @(244,275) /sn:0 /w:[ 0 ]
  //: input g9 (A0) @(240,211) /sn:0 /w:[ 0 ]
  //: output g12 (C0) @(512,277) /sn:0 /w:[ 0 ]
  //: output g11 (S0) @(510,224) /sn:0 /w:[ 0 ]

endmodule

module HalfAdder(B, A, S, C);
//: interface  /sz:(183, 127) /bd:[ Li0>A(28/127) Li1>B(91/127) Ro0<S(39/127) Ro1<C(93/127) ]
input B;    //: /sn:0 {0}(10,58)(21,58){1}
//: {2}(25,58)(45,58)(45,49)(53,49){3}
//: {4}(23,60)(23,80)(54,80){5}
input A;    //: /sn:0 {0}(10,44)(31,44){1}
//: {2}(35,44)(53,44){3}
//: {4}(33,46)(33,75)(54,75){5}
output C;    //: /sn:0 {0}(75,78)(100,78){1}
output S;    //: /sn:0 {0}(99,47)(74,47){1}
//: enddecls

  //: joint g4 (A) @(33, 44) /w:[ 2 -1 1 4 ]
  //: input g3 (B) @(8,58) /sn:0 /w:[ 0 ]
  //: input g2 (A) @(8,44) /sn:0 /w:[ 0 ]
  xor g1 (.I0(A), .I1(B), .Z(S));   //: @(64,47) /sn:0 /delay:" 2" /w:[ 3 3 1 ]
  //: output g6 (S) @(96,47) /sn:0 /w:[ 0 ]
  //: output g7 (C) @(97,78) /sn:0 /w:[ 1 ]
  //: joint g5 (B) @(23, 58) /w:[ 2 -1 1 4 ]
  and g0 (.I0(A), .I1(B), .Z(C));   //: @(65,78) /sn:0 /w:[ 5 5 0 ]

endmodule
