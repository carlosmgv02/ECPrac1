//: version "1.8.7"

module ha(S, CO, B, A);
//: interface  /sz:(55, 65) /bd:[ Li0>A(20/65) Li1>B(35/65) Ro0<S(21/65) Ro1<CO(41/65) ]
input B;    //: /sn:0 {0}(170,290)(233,290)(233,291)(292,291){1}
//: {2}(296,291)(373,291)(373,258)(377,258){3}
//: {4}(294,289)(294,259)(302,259){5}
input A;    //: /sn:0 {0}(171,218)(275,218){1}
//: {2}(279,218)(365,218)(365,253)(377,253){3}
//: {4}(277,220)(277,254)(302,254){5}
output CO;    //: /sn:0 /dp:1 {0}(323,257)(352,257){1}
output S;    //: /sn:0 {0}(428,255)(407,255)(407,256)(398,256){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(388,256) /sn:0 /delay:" 2" /w:[ 3 3 1 ]
  //: output g3 (S) @(425,255) /sn:0 /w:[ 0 ]
  //: output g2 (CO) @(349,257) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(168,290) /sn:0 /w:[ 0 ]
  //: joint g6 (A) @(277, 218) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(294, 291) /w:[ 2 4 1 -1 ]
  and g5 (.I0(A), .I1(B), .Z(CO));   //: @(313,257) /sn:0 /tech:unit /w:[ 5 5 0 ]
  //: input g0 (A) @(169,218) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire w4;    //: /sn:0 {0}(59,96)(96,96){1}
wire w3;    //: /sn:0 {0}(153,126)(235,126)(235,88){1}
wire w2;    //: /sn:0 {0}(153,94)(202,94)(202,80){1}
wire w5;    //: /sn:0 {0}(60,125)(96,125){1}
//: enddecls

  //: switch g4 (w5) @(43,125) /sn:0 /w:[ 0 ] /st:1
  //: switch g3 (w4) @(42,96) /sn:0 /w:[ 0 ] /st:1
  led g2 (.I(w3));   //: @(235,81) /sn:0 /w:[ 1 ] /type:0
  led g1 (.I(w2));   //: @(202,73) /sn:0 /w:[ 1 ] /type:0
  ha g0 (.B(w5), .A(w4), .CO(w3), .S(w2));   //: @(97, 78) /sz:(55, 65) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]

endmodule
