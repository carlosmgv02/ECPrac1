//: version "1.8.7"

module main;    //: root_module
wire w6;    //: /sn:0 {0}(79,61)(107,61)(107,90){1}
wire w4;    //: /sn:0 {0}(113,168)(113,223)(133,223)(133,213){1}
wire w3;    //: /sn:0 {0}(183,168)(183,228)(210,228)(210,218){1}
wire w0;    //: /sn:0 {0}(140,26)(178,26)(178,90){1}
wire w1;    //: /sn:0 {0}(253,68)(263,68)(263,120)(220,120){1}
wire w5;    //: /sn:0 {0}(147,168)(147,224)(167,224)(167,214){1}
//: enddecls

  led g4 (.I(w4));   //: @(133,206) /sn:0 /w:[ 1 ] /type:0
  //: switch g3 (w1) @(236,68) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w0) @(123,26) /sn:0 /w:[ 0 ] /st:0
  //: switch g1 (w6) @(62,61) /sn:0 /w:[ 0 ] /st:0
  led g6 (.I(w3));   //: @(210,211) /sn:0 /w:[ 1 ] /type:0
  led g5 (.I(w5));   //: @(167,207) /sn:0 /w:[ 1 ] /type:0
  PFA_v2 g0 (.B(w0), .A(w6), .C(w1), .G(w5), .P(w4), .S(w3));   //: @(85, 91) /sz:(134, 76) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Bo0<0 Bo1<0 Bo2<0 ]

endmodule

module PFA(C, B, G, S, P, A);
//: interface  /sz:(134, 76) /bd:[ Ti0>A(22/134) Ti1>B(93/134) Ri0>C(29/76) Bo0<S(98/134) Bo1<P(28/134) Bo2<G(62/134) ]
input B;    //: /sn:0 {0}(79,146)(105,146){1}
//: {2}(109,146)(156,146)(156,108)(164,108){3}
//: {4}(107,148)(107,261)(181,261){5}
input A;    //: /sn:0 {0}(88,93)(134,93){1}
//: {2}(138,93)(156,93)(156,103)(164,103){3}
//: {4}(136,95)(136,256)(181,256){5}
output G;    //: /sn:0 /dp:1 {0}(202,259)(268,259)(268,256)(278,256){1}
output P;    //: /sn:0 /dp:1 {0}(185,106)(216,106)(216,94)(220,94){1}
//: {2}(224,94)(229,94)(229,112)(232,112){3}
//: {4}(222,92)(222,71)(293,71){5}
input C;    //: /sn:0 {0}(91,219)(222,219)(222,117)(232,117){1}
output S;    //: /sn:0 /dp:1 {0}(253,115)(297,115){1}
//: enddecls

  and g8 (.I0(A), .I1(B), .Z(G));   //: @(192,259) /sn:0 /delay:" 1" /w:[ 5 5 0 ]
  xor g4 (.I0(P), .I1(C), .Z(S));   //: @(243,115) /sn:0 /delay:" 2" /w:[ 3 1 0 ]
  xor g3 (.I0(A), .I1(B), .Z(P));   //: @(175,106) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  //: input g2 (C) @(89,219) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(77,146) /sn:0 /w:[ 0 ]
  //: output g11 (G) @(275,256) /sn:0 /w:[ 1 ]
  //: joint g10 (B) @(107, 146) /w:[ 2 -1 1 4 ]
  //: joint g6 (P) @(222, 94) /w:[ 2 4 1 -1 ]
  //: joint g9 (A) @(136, 93) /w:[ 2 -1 1 4 ]
  //: output g7 (S) @(294,115) /sn:0 /w:[ 1 ]
  //: output g5 (P) @(290,71) /sn:0 /w:[ 5 ]
  //: input g0 (A) @(86,93) /sn:0 /w:[ 0 ]

endmodule
