//: version "1.8.7"

module HalfAdd(B, A, S, C);
//: interface  /sz:(88, 71) /bd:[ Li0>B(55/71) Li1>A(16/71) Ro0<C(59/71) Ro1<S(12/71) ]
input B;    //: /sn:0 {0}(158,202)(250,202){1}
//: {2}(254,202)(320,202)(320,184)(328,184){3}
//: {4}(252,204)(252,248)(337,248){5}
input A;    //: /sn:0 {0}(157,155)(280,155){1}
//: {2}(284,155)(320,155)(320,179)(328,179){3}
//: {4}(282,157)(282,243)(337,243){5}
output C;    //: /sn:0 {0}(449,246)(358,246){1}
output S;    //: /sn:0 {0}(445,182)(349,182){1}
//: enddecls

  //: joint g4 (A) @(282, 155) /w:[ 2 -1 1 4 ]
  //: input g3 (B) @(156,202) /sn:0 /w:[ 0 ]
  //: input g2 (A) @(155,155) /sn:0 /w:[ 0 ]
  xor g1 (.I0(A), .I1(B), .Z(S));   //: @(339,182) /sn:0 /delay:" 2" /w:[ 3 3 1 ]
  //: output g6 (S) @(442,182) /sn:0 /w:[ 0 ]
  //: output g7 (C) @(446,246) /sn:0 /w:[ 0 ]
  //: joint g5 (B) @(252, 202) /w:[ 2 -1 1 4 ]
  and g0 (.I0(A), .I1(B), .Z(C));   //: @(348,246) /sn:0 /delay:" 1" /w:[ 5 5 1 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 /dp:1 {0}(549,274)(573,274)(573,247){1}
wire w0;    //: /sn:0 {0}(593,121)(593,162){1}
wire w1;    //: /sn:0 {0}(657,205)(614,205){1}
wire w2;    //: /sn:0 /dp:1 {0}(494,186)(494,203)(529,203){1}
wire w5;    //: /sn:0 {0}(549,121)(549,162){1}
//: enddecls

  led g4 (.I(w2));   //: @(494,179) /sn:0 /w:[ 0 ] /type:3
  //: switch g3 (w1) @(675,205) /sn:0 /R:2 /w:[ 0 ] /st:0
  //: switch g2 (w0) @(593,108) /sn:0 /R:3 /w:[ 0 ] /st:1
  //: switch g1 (w5) @(549,108) /sn:0 /R:3 /w:[ 0 ] /st:1
  led g5 (.I(w6));   //: @(542,274) /sn:0 /R:1 /w:[ 0 ] /type:3
  FullAdd g0 (.B(w0), .A(w5), .Cin(w1), .Cout(w2), .S(w6));   //: @(530, 163) /sz:(83, 83) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]

endmodule

module FullAdd(S, Cout, Cin, B, A);
//: interface  /sz:(83, 83) /bd:[ Ti0>B(63/83) Ti1>A(19/83) Ri0>Cin(42/83) Lo0<Cout(40/83) Bo0<S(43/83) ]
input B;    //: /sn:0 {0}(163,178)(214,178)(214,164)(224,164){1}
input A;    //: /sn:0 {0}(161,128)(224,128){1}
output Cout;    //: /sn:0 {0}(606,274)(567,274){1}
input Cin;    //: /sn:0 {0}(394,222)(182,222)(182,246)(165,246){1}
output S;    //: /sn:0 {0}(565,137)(500,137)(500,185)(484,185){1}
wire w3;    //: /sn:0 /dp:1 {0}(546,276)(318,276)(318,168)(308,168){1}
wire w2;    //: /sn:0 /dp:1 {0}(546,271)(494,271)(494,225)(484,225){1}
wire w5;    //: /sn:0 {0}(308,125)(386,125)(386,188)(394,188){1}
//: enddecls

  //: output g4 (S) @(562,137) /sn:0 /w:[ 0 ]
  //: output g3 (Cout) @(603,274) /sn:0 /w:[ 0 ]
  //: input g2 (Cin) @(163,246) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(161,178) /sn:0 /w:[ 0 ]
  HalfAdd g6 (.A(w5), .B(Cin), .S(S), .C(w2));   //: @(395, 174) /sz:(88, 62) /sn:0 /p:[ Li0>1 Li1>0 Ro0<1 Ro1<1 ]
  or g7 (.I0(w2), .I1(w3), .Z(Cout));   //: @(557,274) /sn:0 /w:[ 0 0 1 ]
  HalfAdd g5 (.A(A), .B(B), .S(w5), .C(w3));   //: @(225, 113) /sz:(82, 66) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<1 ]
  //: input g0 (A) @(159,128) /sn:0 /w:[ 0 ]

endmodule
