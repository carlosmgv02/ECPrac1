//: version "1.8.7"

module PFA1(A, Gi, Cin, S, B, Pi);
//: interface  /sz:(68, 63) /bd:[ Ti0>B(52/68) Ti1>A(12/68) Ti2>B(52/68) Ti3>A(12/68) Ri0>Ci(34/63) Ri1>Ci(34/63) Bo0<Gi(9/68) Bo1<Pi(36/68) Bo2<S(57/68) Bo3<Gi(9/68) Bo4<Pi(36/68) Bo5<S(57/68) ]
input B;    //: /sn:0 {0}(120,118)(132,118){1}
//: {2}(136,118)(157,118)(157,102)(166,102){3}
//: {4}(134,120)(134,197){5}
//: {6}(136,199)(194,199)(194,184)(252,184){7}
//: {8}(134,201)(134,242)(257,242){9}
output Gi;    //: /sn:0 {0}(378,240)(278,240){1}
input A;    //: /sn:0 {0}(122,88)(144,88){1}
//: {2}(148,88)(154,88)(154,97)(166,97){3}
//: {4}(146,90)(146,179)(171,179){5}
//: {6}(175,179)(252,179){7}
//: {8}(173,181)(173,237)(257,237){9}
output Pi;    //: /sn:0 {0}(374,182)(273,182){1}
input Cin;    //: /sn:0 {0}(122,152)(254,152)(254,115)(300,115){1}
output S;    //: /sn:0 {0}(394,113)(321,113){1}
wire w3;    //: /sn:0 {0}(300,110)(203,110)(203,100)(187,100){1}
//: enddecls

  //: input g4 (A) @(120,88) /sn:0 /w:[ 0 ]
  //: joint g8 (A) @(146, 88) /w:[ 2 -1 1 4 ]
  and g3 (.I0(A), .I1(B), .Z(Gi));   //: @(268,240) /sn:0 /delay:" 1" /w:[ 9 9 1 ]
  //: output g13 (Gi) @(375,240) /sn:0 /w:[ 0 ]
  or g2 (.I0(A), .I1(B), .Z(Pi));   //: @(263,182) /sn:0 /delay:" 1" /w:[ 7 7 1 ]
  xor g1 (.I0(w3), .I1(Cin), .Z(S));   //: @(311,113) /sn:0 /delay:" 2" /w:[ 0 1 1 ]
  //: joint g11 (B) @(134, 199) /w:[ 6 5 -1 8 ]
  //: joint g10 (B) @(134, 118) /w:[ 2 -1 1 4 ]
  //: input g6 (Cin) @(120,152) /sn:0 /w:[ 0 ]
  //: output g7 (S) @(391,113) /sn:0 /w:[ 0 ]
  //: joint g9 (A) @(173, 179) /w:[ 6 -1 5 8 ]
  //: input g5 (B) @(118,118) /sn:0 /w:[ 0 ]
  xor g0 (.I0(A), .I1(B), .Z(w3));   //: @(177,100) /sn:0 /delay:" 2" /w:[ 3 3 1 ]
  //: output g12 (Pi) @(371,182) /sn:0 /w:[ 0 ]

endmodule

module CLA1(A, C4, S, C0, B);
//: interface  /sz:(168, 40) /bd:[ Ti0>A[3:0](51/168) Ti1>B[3:0](127/168) Ri0>C0(24/40) Lo0<C4(25/40) Bo0<S[3:0](82/168) ]
input [3:0] B;    //: /sn:0 {0}(201,75)(285,75){1}
//: {2}(286,75)(407,75){3}
//: {4}(408,75)(512,75){5}
//: {6}(513,75)(619,75){7}
//: {8}(620,75)(646,75){9}
input C0;    //: /sn:0 {0}(760,176)(690,176)(690,176)(701,176){1}
//: {2}(697,176)(642,176){3}
//: {4}(699,178)(699,276)(662,276){5}
input [3:0] A;    //: /sn:0 {0}(200,55)(251,55){1}
//: {2}(252,55)(367,55){3}
//: {4}(368,55)(471,55){5}
//: {6}(472,55)(586,55){7}
//: {8}(587,55)(643,55){9}
output C4;    //: /sn:0 {0}(167,279)(283,279)(283,279)(232,279){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(817,353)(882,353){1}
wire S1;    //: /sn:0 {0}(811,358)(522,358)(522,206){1}
wire Cin0;    //: /sn:0 {0}(324,255)(324,177)(306,177){1}
wire w16;    //: /sn:0 {0}(501,206)(501,255){1}
wire w15;    //: /sn:0 {0}(368,59)(368,67)(369,67)(369,141){1}
wire w4;    //: /sn:0 {0}(273,207)(273,255){1}
wire w3;    //: /sn:0 {0}(252,59)(252,67)(249,67)(249,143){1}
wire w21;    //: /sn:0 {0}(408,79)(408,87)(409,87)(409,141){1}
wire w28;    //: /sn:0 {0}(587,59)(587,67)(585,67)(585,141){1}
wire w23;    //: /sn:0 {0}(582,206)(582,255){1}
wire S0;    //: /sn:0 {0}(811,368)(630,368)(630,206){1}
wire w22;    //: /sn:0 {0}(609,206)(609,255){1}
wire w17;    //: /sn:0 {0}(478,206)(478,255){1}
wire Cin1;    //: /sn:0 {0}(558,255)(558,176)(534,176){1}
wire w11;    //: /sn:0 {0}(366,206)(366,255){1}
wire Cin;    //: /sn:0 {0}(445,255)(445,176)(426,176){1}
wire w10;    //: /sn:0 {0}(393,206)(393,255){1}
wire w27;    //: /sn:0 {0}(513,79)(513,87)(517,87)(517,141){1}
wire w5;    //: /sn:0 {0}(246,207)(246,255){1}
wire w29;    //: /sn:0 {0}(620,79)(620,87)(625,87)(625,141){1}
wire S3;    //: /sn:0 {0}(811,338)(294,338)(294,207){1}
wire w9;    //: /sn:0 {0}(286,79)(286,87)(289,87)(289,143){1}
wire w26;    //: /sn:0 {0}(472,59)(472,67)(477,67)(477,141){1}
wire S2;    //: /sn:0 {0}(811,348)(414,348)(414,206){1}
//: enddecls

  concat g8 (.I0(S0), .I1(S1), .I2(S2), .I3(S3), .Z(S));   //: @(816,353) /sn:0 /w:[ 0 0 0 0 0 ] /dr:0
  CLL g4 (.P3(w5), .G3(w4), .P2(w11), .G2(w10), .P1(w17), .G1(w16), .P0(w23), .G0(w22), .C0(C0), .C1(Cin1), .C2(Cin), .C3(Cin0), .C4(C4));   //: @(233, 256) /sz:(428, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>5 To0<0 To1<0 To2<0 Lo0<1 ]
  tran g13(.Z(w3), .I(A[3]));   //: @(252,53) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  PFA1 g3 (.B(w29), .A(w28), .Cin(C0), .Gi(w23), .Pi(w22), .S(S0));   //: @(573, 142) /sz:(68, 63) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>3 Bo0<0 Bo1<0 Bo2<1 ]
  PFA1 g2 (.B(w27), .A(w26), .Cin(Cin1), .Gi(w17), .Pi(w16), .S(S1));   //: @(465, 142) /sz:(68, 63) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Bo0<0 Bo1<0 Bo2<1 ]
  PFA1 g1 (.B(w21), .A(w15), .Cin(Cin), .Gi(w11), .Pi(w10), .S(S2));   //: @(357, 142) /sz:(68, 63) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Bo0<0 Bo1<0 Bo2<1 ]
  tran g16(.Z(w21), .I(B[2]));   //: @(408,73) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: input g11 (A) @(198,55) /sn:0 /w:[ 0 ]
  //: output g6 (C4) @(170,279) /sn:0 /R:2 /w:[ 0 ]
  //: joint g9 (C0) @(699, 176) /w:[ 1 -1 2 4 ]
  //: output g7 (S) @(879,353) /sn:0 /w:[ 1 ]
  tran g20(.Z(w28), .I(A[0]));   //: @(587,53) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g15(.Z(w15), .I(A[2]));   //: @(368,53) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g17(.Z(w26), .I(A[1]));   //: @(472,53) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: input g5 (C0) @(762,176) /sn:0 /R:2 /w:[ 0 ]
  tran g14(.Z(w9), .I(B[3]));   //: @(286,73) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g21(.Z(w29), .I(B[0]));   //: @(620,73) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  PFA1 g0 (.B(w9), .A(w3), .Cin(Cin0), .Gi(w5), .Pi(w4), .S(S3));   //: @(237, 144) /sz:(68, 62) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Bo0<0 Bo1<0 Bo2<1 ]
  tran g18(.Z(w27), .I(B[1]));   //: @(513,73) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: input g12 (B) @(199,75) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire w3;    //: /sn:0 {0}(404,102)(431,102){1}
wire [3:0] w0;    //: /sn:0 {0}(514,154)(514,118){1}
wire [3:0] A;    //: /sn:0 /dp:1 {0}(458,14)(458,65)(483,65)(483,76){1}
wire [3:0] w1;    //: /sn:0 {0}(576,11)(576,65)(559,65)(559,76){1}
wire w2;    //: /sn:0 {0}(636,101)(601,101){1}
//: enddecls

  //: dip B (w1) @(576,1) /sn:0 /w:[ 0 ] /st:0
  led g3 (.I(w0));   //: @(514,161) /sn:0 /R:2 /w:[ 0 ] /type:3
  led g2 (.I(w3));   //: @(397,102) /sn:0 /R:1 /w:[ 0 ] /type:3
  //: switch g1 (w2) @(654,101) /sn:0 /R:2 /w:[ 0 ] /st:1
  //: dip A (A) @(458,4) /sn:0 /w:[ 0 ] /st:1
  CLA1 g0 (.B(w1), .A(A), .C0(w2), .C4(w3), .S(w0));   //: @(432, 77) /sz:(168, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]

endmodule

module CLL(G0, P0, P2, G3, P1, G1, P3, C2, G2, C1, C0, C4, C3);
//: interface  /sz:(428, 40) /bd:[ Ti0>P3(13/428) Ti1>G3(41/428) Ti2>P2(132/428) Ti3>G2(160/428) Ti4>P1(245/428) Ti5>G1(269/428) Ti6>P0(349/428) Ti7>G0(376/428) Ri0>C0(20/40) To0<C1(325/428) To1<C2(212/428) To2<C3(91/428) Lo0<C4(23/40) ]
input G2;    //: /sn:0 {0}(76,339)(153,339){1}
//: {2}(157,339)(341,339)(341,308)(388,308){3}
//: {4}(155,341)(155,454)(240,454){5}
input C0;    //: /sn:0 {0}(78,72)(137,72){1}
//: {2}(141,72)(281,72)(281,90)(289,90){3}
//: {4}(139,74)(139,180)(213,180){5}
//: {6}(217,180)(232,180){7}
//: {8}(215,182)(215,264)(230,264){9}
//: {10}(234,264)(239,264){11}
//: {12}(232,266)(232,353)(241,353){13}
input P1;    //: /sn:0 {0}(241,363)(215,363){1}
//: {2}(211,363)(199,363)(199,300){3}
//: {4}(201,298)(239,298){5}
//: {6}(197,298)(191,298)(191,276){7}
//: {8}(193,274)(239,274){9}
//: {10}(189,274)(148,274)(148,221){11}
//: {12}(150,219)(231,219){13}
//: {14}(146,219)(128,219)(128,192){15}
//: {16}(130,190)(232,190){17}
//: {18}(126,190)(78,190){19}
//: {20}(213,365)(213,398)(242,398){21}
output C3;    //: /sn:0 /dp:1 {0}(409,300)(579,300){1}
input G0;    //: /sn:0 {0}(78,148)(179,148){1}
//: {2}(183,148)(324,148)(324,107)(408,107){3}
//: {4}(181,150)(181,214)(202,214){5}
//: {6}(206,214)(231,214){7}
//: {8}(204,216)(204,293)(220,293){9}
//: {10}(224,293)(239,293){11}
//: {12}(222,295)(222,393)(242,393){13}
output C4;    //: /sn:0 /dp:1 {0}(414,402)(589,402){1}
output C2;    //: /sn:0 {0}(576,200)(493,200)(493,201)(408,201){1}
input P3;    //: /sn:0 {0}(241,434)(203,434)(203,410){1}
//: {2}(205,408)(242,408){3}
//: {4}(201,408)(187,408)(187,375){5}
//: {6}(189,373)(241,373){7}
//: {8}(185,373)(76,373){9}
input G1;    //: /sn:0 {0}(77,239)(138,239){1}
//: {2}(142,239)(290,239)(290,206)(387,206){3}
//: {4}(140,241)(140,321)(167,321){5}
//: {6}(171,321)(205,321)(205,321)(239,321){7}
//: {8}(169,323)(169,424)(241,424){9}
input G3;    //: /sn:0 {0}(78,436)(118,436)(118,459)(240,459){1}
input P0;    //: /sn:0 {0}(78,111)(97,111){1}
//: {2}(101,111)(281,111)(281,95)(289,95){3}
//: {4}(99,113)(99,185)(159,185){5}
//: {6}(163,185)(232,185){7}
//: {8}(161,187)(161,269)(208,269){9}
//: {10}(212,269)(239,269){11}
//: {12}(210,271)(210,358)(241,358){13}
output C1;    //: /sn:0 {0}(572,105)(429,105){1}
input P2;    //: /sn:0 {0}(242,403)(222,403){1}
//: {2}(218,403)(205,403)(205,370){3}
//: {4}(207,368)(241,368){5}
//: {6}(203,368)(191,368)(191,328){7}
//: {8}(193,326)(216,326)(216,326)(239,326){9}
//: {10}(189,326)(185,326)(185,305){11}
//: {12}(187,303)(239,303){13}
//: {14}(183,303)(175,303)(175,281){15}
//: {16}(177,279)(239,279){17}
//: {18}(173,279)(78,279){19}
//: {20}(220,405)(220,429)(241,429){21}
wire w6;    //: /sn:0 /dp:1 {0}(393,400)(263,400){1}
wire w7;    //: /sn:0 {0}(262,363)(383,363)(383,395)(393,395){1}
wire w14;    //: /sn:0 {0}(393,410)(357,410)(357,457)(261,457){1}
wire w4;    //: /sn:0 /dp:1 {0}(388,298)(260,298){1}
wire w3;    //: /sn:0 {0}(253,185)(377,185)(377,196)(387,196){1}
wire w1;    //: /sn:0 /dp:1 {0}(387,201)(265,201)(265,217)(252,217){1}
wire w2;    //: /sn:0 {0}(310,93)(398,93)(398,102)(408,102){1}
wire w10;    //: /sn:0 {0}(262,429)(327,429)(327,405)(393,405){1}
wire w5;    //: /sn:0 {0}(260,271)(378,271)(378,293)(388,293){1}
wire w9;    //: /sn:0 {0}(388,303)(323,303)(323,324)(260,324){1}
//: enddecls

  or g4 (.I0(w2), .I1(G0), .Z(C1));   //: @(419,105) /sn:0 /delay:" 1" /w:[ 1 3 1 ]
  and g8 (.I0(C0), .I1(P0), .I2(P1), .Z(w3));   //: @(243,185) /sn:0 /delay:" 1" /w:[ 7 7 17 0 ]
  //: joint g37 (P1) @(199, 298) /w:[ 4 -1 6 3 ]
  and g34 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .I4(P3), .Z(w7));   //: @(252,363) /sn:0 /delay:" 1" /w:[ 13 13 0 5 7 0 ]
  and g3 (.I0(C0), .I1(P0), .Z(w2));   //: @(300,93) /sn:0 /delay:" 1" /w:[ 3 3 0 ]
  //: joint g13 (G0) @(181, 148) /w:[ 2 -1 1 4 ]
  //: input g2 (G0) @(76,148) /sn:0 /w:[ 0 ]
  //: input g1 (P0) @(76,111) /sn:0 /w:[ 0 ]
  and g11 (.I0(G0), .I1(P1), .Z(w1));   //: @(242,217) /sn:0 /delay:" 1" /w:[ 7 13 1 ]
  //: input g16 (P2) @(76,279) /sn:0 /w:[ 19 ]
  or g50 (.I0(w7), .I1(w6), .I2(w10), .I3(w14), .Z(C4));   //: @(404,402) /sn:0 /delay:" 1" /w:[ 1 0 1 0 0 ]
  //: joint g28 (P2) @(185, 303) /w:[ 12 -1 14 11 ]
  //: joint g10 (C0) @(139, 72) /w:[ 2 -1 1 4 ]
  //: input g32 (G3) @(76,436) /sn:0 /w:[ 0 ]
  //: joint g27 (G1) @(140, 239) /w:[ 2 -1 1 4 ]
  //: joint g19 (C0) @(215, 180) /w:[ 6 -1 5 8 ]
  //: joint g38 (P2) @(191, 326) /w:[ 8 -1 10 7 ]
  //: input g6 (P1) @(76,190) /sn:0 /w:[ 19 ]
  //: input g7 (G1) @(75,239) /sn:0 /w:[ 0 ]
  //: joint g9 (P0) @(99, 111) /w:[ 2 -1 1 4 ]
  //: input g31 (P3) @(74,373) /sn:0 /w:[ 9 ]
  //: joint g20 (P0) @(161, 185) /w:[ 6 -1 5 8 ]
  //: output g15 (C2) @(573,200) /sn:0 /w:[ 0 ]
  and g39 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w6));   //: @(253,400) /sn:0 /delay:" 1" /w:[ 13 21 0 3 1 ]
  and g48 (.I0(G2), .I1(G3), .Z(w14));   //: @(251,457) /sn:0 /delay:" 1" /w:[ 5 1 1 ]
  //: joint g43 (P3) @(187, 373) /w:[ 6 -1 8 5 ]
  or g29 (.I0(w5), .I1(w4), .I2(w9), .I3(G2), .Z(C3));   //: @(399,300) /sn:0 /delay:" 1" /w:[ 1 0 0 3 0 ]
  //: joint g25 (P2) @(175, 279) /w:[ 16 -1 18 15 ]
  //: input g17 (G2) @(74,339) /sn:0 /w:[ 0 ]
  //: joint g42 (P2) @(205, 368) /w:[ 4 -1 6 3 ]
  //: output g5 (C1) @(569,105) /sn:0 /w:[ 0 ]
  or g14 (.I0(w3), .I1(w1), .I2(G1), .Z(C2));   //: @(398,201) /sn:0 /delay:" 1" /w:[ 1 0 3 1 ]
  //: joint g47 (P3) @(203, 408) /w:[ 2 -1 4 1 ]
  and g44 (.I0(G1), .I1(P2), .I2(P3), .Z(w10));   //: @(252,429) /sn:0 /delay:" 1" /w:[ 9 21 0 0 ]
  //: joint g36 (P0) @(210, 269) /w:[ 10 -1 9 12 ]
  //: joint g24 (P1) @(191, 274) /w:[ 8 -1 10 7 ]
  //: joint g21 (P1) @(148, 219) /w:[ 12 -1 14 11 ]
  //: joint g41 (P1) @(213, 363) /w:[ 1 -1 2 20 ]
  //: joint g23 (G0) @(204, 214) /w:[ 6 -1 5 8 ]
  //: joint g40 (G0) @(222, 293) /w:[ 10 -1 9 12 ]
  //: joint g46 (P2) @(220, 403) /w:[ 1 -1 2 20 ]
  //: joint g45 (G1) @(169, 321) /w:[ 6 -1 5 8 ]
  //: joint g35 (C0) @(232, 264) /w:[ 10 -1 9 12 ]
  and g26 (.I0(G1), .I1(P2), .Z(w9));   //: @(250,324) /sn:0 /delay:" 1" /w:[ 7 9 1 ]
  and g22 (.I0(G0), .I1(P1), .I2(P2), .Z(w4));   //: @(250,298) /sn:0 /delay:" 1" /w:[ 11 5 13 1 ]
  //: input g0 (C0) @(76,72) /sn:0 /w:[ 0 ]
  //: joint g12 (P1) @(128, 190) /w:[ 16 -1 18 15 ]
  and g18 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .Z(w5));   //: @(250,271) /sn:0 /delay:" 1" /w:[ 11 11 9 17 0 ]
  //: output g33 (C4) @(586,402) /sn:0 /w:[ 1 ]
  //: output g30 (C3) @(576,300) /sn:0 /w:[ 1 ]
  //: joint g49 (G2) @(155, 339) /w:[ 2 -1 1 4 ]

endmodule
