//: version "1.8.7"

module PFA1(A, Gi, Cin, S, B, Pi);
//: interface  /sz:(68, 63) /bd:[ Ti0>A(12/68) Ti1>B(52/68) Ri0>Ci(34/63) Bo0<S(57/68) Bo1<Pi(36/68) Bo2<Gi(9/68) ]
input B;    //: /sn:0 {0}(120,118)(132,118){1}
//: {2}(136,118)(157,118)(157,102)(166,102){3}
//: {4}(134,120)(134,197){5}
//: {6}(136,199)(194,199)(194,184)(252,184){7}
//: {8}(134,201)(134,242)(257,242){9}
output Gi;    //: /sn:0 {0}(378,240)(278,240){1}
input A;    //: /sn:0 {0}(122,88)(144,88){1}
//: {2}(148,88)(154,88)(154,97)(166,97){3}
//: {4}(146,90)(146,179)(171,179){5}
//: {6}(175,179)(252,179){7}
//: {8}(173,181)(173,237)(257,237){9}
output Pi;    //: /sn:0 {0}(374,182)(273,182){1}
input Cin;    //: /sn:0 {0}(122,152)(253,152)(253,115)(300,115){1}
output S;    //: /sn:0 {0}(394,113)(321,113){1}
wire w3;    //: /sn:0 {0}(300,110)(203,110)(203,100)(187,100){1}
//: enddecls

  //: joint g8 (A) @(146, 88) /w:[ 2 -1 1 4 ]
  //: input g4 (A) @(120,88) /sn:0 /w:[ 0 ]
  //: output g13 (Gi) @(375,240) /sn:0 /w:[ 0 ]
  and g3 (.I0(A), .I1(B), .Z(Gi));   //: @(268,240) /sn:0 /delay:" 1" /w:[ 9 9 1 ]
  or g2 (.I0(A), .I1(B), .Z(Pi));   //: @(263,182) /sn:0 /delay:" 1" /w:[ 7 7 1 ]
  xor g1 (.I0(w3), .I1(Cin), .Z(S));   //: @(311,113) /sn:0 /delay:" 2" /w:[ 0 1 1 ]
  //: joint g11 (B) @(134, 199) /w:[ 6 5 -1 8 ]
  //: joint g10 (B) @(134, 118) /w:[ 2 -1 1 4 ]
  //: input g6 (Cin) @(120,152) /sn:0 /w:[ 0 ]
  //: joint g9 (A) @(173, 179) /w:[ 6 -1 5 8 ]
  //: output g7 (S) @(391,113) /sn:0 /w:[ 0 ]
  //: input g5 (B) @(118,118) /sn:0 /w:[ 0 ]
  xor g0 (.I0(A), .I1(B), .Z(w3));   //: @(177,100) /sn:0 /delay:" 2" /w:[ 3 3 1 ]
  //: output g12 (Pi) @(371,182) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire B;    //: /sn:0 /dp:1 {0}(26,66)(46,66)(46,58)(82,58){1}
//: {2}(86,58)(107,58)(107,42)(116,42){3}
//: {4}(84,60)(84,137){5}
//: {6}(86,139)(144,139)(144,124)(202,124){7}
//: {8}(84,141)(84,182)(207,182){9}
wire w3;    //: /sn:0 {0}(250,50)(153,50)(153,40)(137,40){1}
wire A;    //: /sn:0 /dp:1 {0}(26,29)(93,29){1}
//: {2}(97,29)(103,29)(103,37)(116,37){3}
//: {4}(95,31)(95,119)(121,119){5}
//: {6}(125,119)(202,119){7}
//: {8}(123,121)(123,177)(207,177){9}
wire w0;    //: /sn:0 {0}(345,53)(271,53){1}
wire w1;    //: /sn:0 {0}(344,122)(223,122){1}
wire w2;    //: /sn:0 {0}(344,180)(228,180){1}
wire Cin;    //: /sn:0 {0}(26,106)(49,106)(49,92)(157,92)(157,55)(250,55){1}
//: enddecls

  //: joint g8 (A) @(95, 29) /w:[ 2 -1 1 4 ]
  led g4 (.I(w0));   //: @(352,53) /sn:0 /R:3 /w:[ 0 ] /type:3
  and g3 (.I0(A), .I1(B), .Z(w2));   //: @(218,180) /sn:0 /delay:" 1" /w:[ 9 9 1 ]
  led g13 (.I(w2));   //: @(351,180) /sn:0 /R:3 /w:[ 0 ] /type:3
  or g2 (.I0(A), .I1(B), .Z(w1));   //: @(213,122) /sn:0 /delay:" 1" /w:[ 7 7 1 ]
  xor g1 (.I0(w3), .I1(Cin), .Z(w0));   //: @(261,53) /sn:0 /delay:" 2" /w:[ 0 1 1 ]
  //: joint g11 (B) @(84, 139) /w:[ 6 5 -1 8 ]
  //: joint g10 (B) @(84, 58) /w:[ 2 -1 1 4 ]
  //: switch g6 (B) @(9,66) /sn:0 /w:[ 0 ] /st:0
  //: joint g9 (A) @(123, 119) /w:[ 6 -1 5 8 ]
  //: switch g7 (Cin) @(9,106) /sn:0 /w:[ 0 ] /st:0
  //: switch g5 (A) @(9,29) /sn:0 /w:[ 0 ] /st:0
  xor g0 (.I0(A), .I1(B), .Z(w3));   //: @(127,40) /sn:0 /delay:" 2" /w:[ 3 3 1 ]
  led g12 (.I(w1));   //: @(351,122) /sn:0 /R:3 /w:[ 0 ] /type:3

endmodule
