//: version "1.8.7"

module PFA2(Si, Ci, Bi, Gi, Pi, Ai);
//: interface  /sz:(75, 67) /bd:[ Ti0>A(20/75) Ti1>B(57/75) Ri0>Ci(35/67) Bo0<Gi(12/75) Bo1<Pi(38/75) Bo2<S(61/75) ]
output Gi;    //: /sn:0 {0}(482,170)(374,170){1}
input Bi;    //: /sn:0 /dp:1 {0}(327,90)(300,90)(300,112)(251,112){1}
//: {2}(247,112)(214,112){3}
//: {4}(249,114)(249,172)(353,172){5}
input Ai;    //: /sn:0 {0}(214,70)(274,70){1}
//: {2}(278,70)(298,70)(298,85)(327,85){3}
//: {4}(276,72)(276,167)(353,167){5}
output Si;    //: /sn:0 {0}(479,117)(423,117){1}
output Pi;    //: /sn:0 {0}(478,88)(377,88){1}
//: {2}(373,88)(348,88){3}
//: {4}(375,90)(375,114)(402,114){5}
input Ci;    //: /sn:0 {0}(216,157)(313,157)(313,119)(402,119){1}
//: enddecls

  xor g4 (.I0(Pi), .I1(Ci), .Z(Si));   //: @(413,117) /sn:0 /delay:" 2" /w:[ 5 1 1 ]
  //: output g8 (Si) @(476,117) /sn:0 /w:[ 0 ]
  xor g3 (.I0(Ai), .I1(Bi), .Z(Pi));   //: @(338,88) /sn:0 /delay:" 2" /w:[ 3 0 3 ]
  //: input g2 (Ci) @(214,157) /sn:0 /w:[ 0 ]
  //: input g1 (Bi) @(212,112) /sn:0 /w:[ 3 ]
  //: output g11 (Gi) @(479,170) /sn:0 /w:[ 0 ]
  //: joint g10 (Bi) @(249, 112) /w:[ 1 -1 2 4 ]
  //: output g6 (Pi) @(475,88) /sn:0 /w:[ 0 ]
  //: joint g7 (Pi) @(375, 88) /w:[ 1 -1 2 4 ]
  //: joint g9 (Ai) @(276, 70) /w:[ 2 -1 1 4 ]
  and g5 (.I0(Ai), .I1(Bi), .Z(Gi));   //: @(364,170) /sn:0 /delay:" 1" /w:[ 5 5 1 ]
  //: input g0 (Ai) @(212,70) /sn:0 /w:[ 0 ]

endmodule

module CLA2(C4, B, A, S, C1);
//: interface  /sz:(243, 46) /bd:[ Ti0>A[3:0](63/243) Ti1>B[3:0](174/243) Ri0>C1(28/46) Lo0<C4(25/46) Bo0<S[3:0](116/243) ]
input [3:0] B;    //: /sn:0 {0}(109,68)(247,68){1}
//: {2}(248,68)(400,68){3}
//: {4}(401,68)(564,68){5}
//: {6}(565,68)(730,68){7}
//: {8}(731,68)(768,68){9}
input [3:0] A;    //: /sn:0 {0}(111,40)(210,40){1}
//: {2}(211,40)(359,40){3}
//: {4}(360,40)(531,40){5}
//: {6}(532,40)(691,40){7}
//: {8}(692,40)(767,40){9}
output C4;    //: /sn:0 {0}(133,300)(174,300){1}
input C1;    //: /sn:0 {0}(828,176)(809,176){1}
//: {2}(805,176)(749,176){3}
//: {4}(807,178)(807,302)(754,302){5}
output [3:0] S;    //: /sn:0 /dp:1 {0}(773,382)(820,382){1}
wire A0;    //: /sn:0 {0}(692,44)(692,52)(693,52)(693,140){1}
wire S1;    //: /sn:0 /dp:1 {0}(569,213)(569,387)(767,387){1}
wire Gi;    //: /sn:0 {0}(685,209)(685,274){1}
wire w16;    //: /sn:0 {0}(228,214)(228,274){1}
wire w14;    //: /sn:0 {0}(265,181)(300,181)(300,274){1}
wire w4;    //: /sn:0 {0}(546,213)(546,274){1}
wire A3;    //: /sn:0 {0}(211,44)(211,52)(209,52)(209,145){1}
wire w0;    //: /sn:0 {0}(250,214)(250,367)(767,367){1}
wire A2;    //: /sn:0 {0}(360,44)(360,52)(365,52)(365,139){1}
wire B2;    //: /sn:0 {0}(401,72)(401,80)(402,80)(402,139){1}
wire w28;    //: /sn:0 {0}(470,274)(470,175)(421,175){1}
wire B1;    //: /sn:0 {0}(565,72)(565,144){1}
wire S0;    //: /sn:0 /dp:1 {0}(734,209)(734,397)(767,397){1}
wire w17;    //: /sn:0 {0}(201,214)(201,274){1}
wire Pi;    //: /sn:0 {0}(711,209)(711,274){1}
wire w11;    //: /sn:0 {0}(357,208)(357,274){1}
wire w2;    //: /sn:0 {0}(584,180)(634,180)(634,274){1}
wire w10;    //: /sn:0 {0}(383,208)(383,274){1}
wire A1;    //: /sn:0 {0}(532,44)(532,52)(528,52)(528,144){1}
wire w5;    //: /sn:0 {0}(520,213)(520,274){1}
wire B3;    //: /sn:0 {0}(248,72)(248,80)(246,80)(246,145){1}
wire B0;    //: /sn:0 {0}(731,72)(731,80)(730,80)(730,140){1}
wire S2;    //: /sn:0 /dp:1 {0}(406,208)(406,377)(767,377){1}
//: enddecls

  CLL g4 (.G3(w17), .P3(w16), .G2(w11), .P2(w10), .P1(w4), .G1(w5), .G0(Gi), .P0(Pi), .C0(C1), .C3(w14), .C2(w28), .C1(w2), .C4(C4));   //: @(175, 275) /sz:(578, 50) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>5 To0<1 To1<0 To2<1 Lo0<1 ]
  PFA2 g3 (.Ai(A3), .Bi(B3), .Ci(w14), .Gi(w17), .Pi(w16), .Si(w0));   //: @(189, 146) /sz:(75, 67) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<0 Bo1<0 Bo2<0 ]
  PFA2 g2 (.Ai(A2), .Bi(B2), .Ci(w28), .Gi(w11), .Pi(w10), .Si(S2));   //: @(345, 140) /sz:(75, 67) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Bo0<0 Bo1<0 Bo2<0 ]
  PFA2 g1 (.Ai(A1), .Bi(B1), .Ci(w2), .Gi(w5), .Pi(w4), .Si(S1));   //: @(508, 145) /sz:(75, 67) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<0 Bo1<0 Bo2<0 ]
  tran g11(.Z(A1), .I(A[1]));   //: @(532,38) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g10(.Z(A2), .I(A[2]));   //: @(360,38) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: output g19 (C4) @(136,300) /sn:0 /R:2 /w:[ 0 ]
  //: joint g6 (C1) @(807, 176) /w:[ 1 -1 2 4 ]
  //: input g7 (B) @(107,68) /sn:0 /w:[ 0 ]
  tran g9(.Z(A3), .I(A[3]));   //: @(211,38) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g15(.Z(B2), .I(B[2]));   //: @(401,66) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g20(.Z(B3), .I(B[3]));   //: @(248,66) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g17(.Z(B1), .I(B[1]));   //: @(565,66) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: input g5 (A) @(109,40) /sn:0 /w:[ 0 ]
  tran g14(.Z(B0), .I(B[0]));   //: @(731,66) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: output g21 (S) @(817,382) /sn:0 /w:[ 1 ]
  concat g23 (.I0(S0), .I1(S1), .I2(S2), .I3(w0), .Z(S));   //: @(772,382) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0
  PFA2 g0 (.Ai(A0), .Bi(B0), .Ci(C1), .Gi(Gi), .Pi(Pi), .Si(S0));   //: @(673, 141) /sz:(75, 67) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>3 Bo0<0 Bo1<0 Bo2<0 ]
  //: input g22 (C1) @(830,176) /sn:0 /R:2 /w:[ 0 ]
  tran g12(.Z(A0), .I(A[0]));   //: @(692,38) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1

endmodule

module main;    //: root_module
wire w4;    //: /sn:0 {0}(218,90)(261,90){1}
wire [3:0] w3;    //: /sn:0 {0}(378,136)(378,112){1}
wire [3:0] w0;    //: /sn:0 /dp:1 {0}(325,26)(325,64){1}
wire [3:0] w1;    //: /sn:0 /dp:1 {0}(436,25)(436,64){1}
wire w2;    //: /sn:0 {0}(558,93)(506,93){1}
//: enddecls

  led g4 (.I(w3));   //: @(378,143) /sn:0 /R:2 /w:[ 0 ] /type:3
  //: switch g3 (w2) @(576,93) /sn:0 /R:2 /w:[ 0 ] /st:1
  //: dip g2 (w1) @(436,15) /sn:0 /w:[ 0 ] /st:0
  //: dip g1 (w0) @(325,16) /sn:0 /w:[ 0 ] /st:0
  led g5 (.I(w4));   //: @(211,90) /sn:0 /R:1 /w:[ 0 ] /type:3
  CLA2 g0 (.B(w1), .A(w0), .C1(w2), .C4(w4), .S(w3));   //: @(262, 65) /sz:(243, 46) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]

endmodule

module CLL(G0, P0, P2, G3, P1, G1, P3, C2, G2, C1, C0, C4, C3);
//: interface  /sz:(40, 40) /bd:[ ]
input G2;    //: /sn:0 {0}(76,339)(153,339){1}
//: {2}(157,339)(341,339)(341,308)(388,308){3}
//: {4}(155,341)(155,454)(240,454){5}
input C0;    //: /sn:0 {0}(78,72)(137,72){1}
//: {2}(141,72)(281,72)(281,90)(289,90){3}
//: {4}(139,74)(139,180)(213,180){5}
//: {6}(217,180)(232,180){7}
//: {8}(215,182)(215,264)(230,264){9}
//: {10}(234,264)(239,264){11}
//: {12}(232,266)(232,353)(241,353){13}
input P1;    //: /sn:0 {0}(241,363)(215,363){1}
//: {2}(211,363)(199,363)(199,300){3}
//: {4}(201,298)(239,298){5}
//: {6}(197,298)(191,298)(191,276){7}
//: {8}(193,274)(239,274){9}
//: {10}(189,274)(148,274)(148,221){11}
//: {12}(150,219)(231,219){13}
//: {14}(146,219)(128,219)(128,192){15}
//: {16}(130,190)(232,190){17}
//: {18}(126,190)(78,190){19}
//: {20}(213,365)(213,398)(242,398){21}
output C3;    //: /sn:0 /dp:1 {0}(409,300)(579,300){1}
input G0;    //: /sn:0 {0}(78,148)(179,148){1}
//: {2}(183,148)(324,148)(324,107)(408,107){3}
//: {4}(181,150)(181,214)(202,214){5}
//: {6}(206,214)(231,214){7}
//: {8}(204,216)(204,293)(220,293){9}
//: {10}(224,293)(239,293){11}
//: {12}(222,295)(222,393)(242,393){13}
output C4;    //: /sn:0 /dp:1 {0}(414,402)(589,402){1}
output C2;    //: /sn:0 {0}(576,200)(493,200)(493,201)(408,201){1}
input P3;    //: /sn:0 {0}(241,434)(203,434)(203,410){1}
//: {2}(205,408)(242,408){3}
//: {4}(201,408)(187,408)(187,375){5}
//: {6}(189,373)(241,373){7}
//: {8}(185,373)(76,373){9}
input G1;    //: /sn:0 {0}(77,239)(138,239){1}
//: {2}(142,239)(290,239)(290,206)(387,206){3}
//: {4}(140,241)(140,321)(167,321){5}
//: {6}(171,321)(205,321)(205,321)(239,321){7}
//: {8}(169,323)(169,424)(241,424){9}
input G3;    //: /sn:0 {0}(78,436)(118,436)(118,459)(240,459){1}
input P0;    //: /sn:0 {0}(78,111)(97,111){1}
//: {2}(101,111)(281,111)(281,95)(289,95){3}
//: {4}(99,113)(99,185)(159,185){5}
//: {6}(163,185)(232,185){7}
//: {8}(161,187)(161,269)(208,269){9}
//: {10}(212,269)(239,269){11}
//: {12}(210,271)(210,358)(241,358){13}
output C1;    //: /sn:0 {0}(572,105)(429,105){1}
input P2;    //: /sn:0 {0}(242,403)(222,403){1}
//: {2}(218,403)(205,403)(205,370){3}
//: {4}(207,368)(241,368){5}
//: {6}(203,368)(191,368)(191,328){7}
//: {8}(193,326)(216,326)(216,326)(239,326){9}
//: {10}(189,326)(185,326)(185,305){11}
//: {12}(187,303)(239,303){13}
//: {14}(183,303)(175,303)(175,281){15}
//: {16}(177,279)(239,279){17}
//: {18}(173,279)(78,279){19}
//: {20}(220,405)(220,429)(241,429){21}
wire w6;    //: /sn:0 /dp:1 {0}(393,400)(263,400){1}
wire w7;    //: /sn:0 {0}(262,363)(383,363)(383,395)(393,395){1}
wire w14;    //: /sn:0 {0}(393,410)(357,410)(357,457)(261,457){1}
wire w4;    //: /sn:0 /dp:1 {0}(388,298)(260,298){1}
wire w3;    //: /sn:0 {0}(253,185)(377,185)(377,196)(387,196){1}
wire w1;    //: /sn:0 /dp:1 {0}(387,201)(265,201)(265,217)(252,217){1}
wire w2;    //: /sn:0 {0}(310,93)(398,93)(398,102)(408,102){1}
wire w10;    //: /sn:0 {0}(262,429)(327,429)(327,405)(393,405){1}
wire w5;    //: /sn:0 {0}(260,271)(378,271)(378,293)(388,293){1}
wire w9;    //: /sn:0 {0}(388,303)(323,303)(323,324)(260,324){1}
//: enddecls

  or g4 (.I0(w2), .I1(G0), .Z(C1));   //: @(419,105) /sn:0 /delay:" 1" /w:[ 1 3 1 ]
  and g8 (.I0(C0), .I1(P0), .I2(P1), .Z(w3));   //: @(243,185) /sn:0 /delay:" 1" /w:[ 7 7 17 0 ]
  //: joint g37 (P1) @(199, 298) /w:[ 4 -1 6 3 ]
  and g34 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .I4(P3), .Z(w7));   //: @(252,363) /sn:0 /delay:" 1" /w:[ 13 13 0 5 7 0 ]
  and g3 (.I0(C0), .I1(P0), .Z(w2));   //: @(300,93) /sn:0 /delay:" 1" /w:[ 3 3 0 ]
  //: joint g13 (G0) @(181, 148) /w:[ 2 -1 1 4 ]
  //: input g2 (G0) @(76,148) /sn:0 /w:[ 0 ]
  //: input g1 (P0) @(76,111) /sn:0 /w:[ 0 ]
  and g11 (.I0(G0), .I1(P1), .Z(w1));   //: @(242,217) /sn:0 /delay:" 1" /w:[ 7 13 1 ]
  //: input g16 (P2) @(76,279) /sn:0 /w:[ 19 ]
  or g50 (.I0(w7), .I1(w6), .I2(w10), .I3(w14), .Z(C4));   //: @(404,402) /sn:0 /delay:" 1" /w:[ 1 0 1 0 0 ]
  //: joint g28 (P2) @(185, 303) /w:[ 12 -1 14 11 ]
  //: joint g10 (C0) @(139, 72) /w:[ 2 -1 1 4 ]
  //: input g32 (G3) @(76,436) /sn:0 /w:[ 0 ]
  //: joint g27 (G1) @(140, 239) /w:[ 2 -1 1 4 ]
  //: joint g19 (C0) @(215, 180) /w:[ 6 -1 5 8 ]
  //: joint g38 (P2) @(191, 326) /w:[ 8 -1 10 7 ]
  //: input g6 (P1) @(76,190) /sn:0 /w:[ 19 ]
  //: input g7 (G1) @(75,239) /sn:0 /w:[ 0 ]
  //: joint g9 (P0) @(99, 111) /w:[ 2 -1 1 4 ]
  //: input g31 (P3) @(74,373) /sn:0 /w:[ 9 ]
  //: joint g20 (P0) @(161, 185) /w:[ 6 -1 5 8 ]
  //: output g15 (C2) @(573,200) /sn:0 /w:[ 0 ]
  and g39 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w6));   //: @(253,400) /sn:0 /delay:" 1" /w:[ 13 21 0 3 1 ]
  and g48 (.I0(G2), .I1(G3), .Z(w14));   //: @(251,457) /sn:0 /delay:" 1" /w:[ 5 1 1 ]
  //: joint g43 (P3) @(187, 373) /w:[ 6 -1 8 5 ]
  or g29 (.I0(w5), .I1(w4), .I2(w9), .I3(G2), .Z(C3));   //: @(399,300) /sn:0 /delay:" 1" /w:[ 1 0 0 3 0 ]
  //: joint g25 (P2) @(175, 279) /w:[ 16 -1 18 15 ]
  //: input g17 (G2) @(74,339) /sn:0 /w:[ 0 ]
  //: joint g42 (P2) @(205, 368) /w:[ 4 -1 6 3 ]
  //: output g5 (C1) @(569,105) /sn:0 /w:[ 0 ]
  or g14 (.I0(w3), .I1(w1), .I2(G1), .Z(C2));   //: @(398,201) /sn:0 /delay:" 1" /w:[ 1 0 3 1 ]
  //: joint g47 (P3) @(203, 408) /w:[ 2 -1 4 1 ]
  and g44 (.I0(G1), .I1(P2), .I2(P3), .Z(w10));   //: @(252,429) /sn:0 /delay:" 1" /w:[ 9 21 0 0 ]
  //: joint g36 (P0) @(210, 269) /w:[ 10 -1 9 12 ]
  //: joint g24 (P1) @(191, 274) /w:[ 8 -1 10 7 ]
  //: joint g21 (P1) @(148, 219) /w:[ 12 -1 14 11 ]
  //: joint g41 (P1) @(213, 363) /w:[ 1 -1 2 20 ]
  //: joint g23 (G0) @(204, 214) /w:[ 6 -1 5 8 ]
  //: joint g40 (G0) @(222, 293) /w:[ 10 -1 9 12 ]
  //: joint g46 (P2) @(220, 403) /w:[ 1 -1 2 20 ]
  //: joint g45 (G1) @(169, 321) /w:[ 6 -1 5 8 ]
  //: joint g35 (C0) @(232, 264) /w:[ 10 -1 9 12 ]
  and g26 (.I0(G1), .I1(P2), .Z(w9));   //: @(250,324) /sn:0 /delay:" 1" /w:[ 7 9 1 ]
  and g22 (.I0(G0), .I1(P1), .I2(P2), .Z(w4));   //: @(250,298) /sn:0 /delay:" 1" /w:[ 11 5 13 1 ]
  //: input g0 (C0) @(76,72) /sn:0 /w:[ 0 ]
  //: joint g12 (P1) @(128, 190) /w:[ 16 -1 18 15 ]
  and g18 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .Z(w5));   //: @(250,271) /sn:0 /delay:" 1" /w:[ 11 11 9 17 0 ]
  //: output g33 (C4) @(586,402) /sn:0 /w:[ 1 ]
  //: output g30 (C3) @(576,300) /sn:0 /w:[ 1 ]
  //: joint g49 (G2) @(155, 339) /w:[ 2 -1 1 4 ]

endmodule
