//: version "1.8.7"
//: property discardChanges = 1

module MAIN();
//: interface  /sz:(40, 40) /bd:[ ]
wire w4;    //: /sn:0 {0}(352,211)(352,179){1}
wire [3:0] w3;    //: /sn:0 {0}(250,211)(250,194)(93,194)(93,108){1}
wire w0;    //: /sn:0 {0}(320,211)(320,191)(333,191)(333,353){1}
wire [3:0] w2;    //: /sn:0 {0}(271,211)(271,181)(183,181)(183,108){1}
wire [3:0] w5;    //: /sn:0 /dp:1 {0}(288,110)(288,182)(289,182)(289,211){1}
//: enddecls

  //: switch g4 (w0) @(333,367) /sn:0 /R:1 /w:[ 1 ] /st:0
  led g3 (.I(w5));   //: @(288,103) /sn:0 /w:[ 0 ] /type:2
  //: dip g2 (w2) @(183,98) /sn:0 /w:[ 1 ] /st:0
  //: dip g1 (w3) @(93,98) /sn:0 /w:[ 1 ] /st:0
  led g5 (.I(w4));   //: @(352,172) /sn:0 /w:[ 1 ] /type:0
  CSA g0 (.A(w3), .B(w2), .Cin(w0), .Cout(w4), .S(w5));   //: @(241, 212) /sz:(127, 64) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 To0<0 To1<1 ]

endmodule

module CSA(B, A, Cin, S, Cout);
//: interface  /sz:(127, 64) /bd:[ Ti0>Cin(74/127) Ti1>B[3:0](30/127) Ti2>A[3:0](9/127) To0<S[3:0](48/127) To1<Cout(96/127) ]
input [3:0] B;    //: /sn:0 /dp:9 {0}(42,44)(143,44){1}
//: {2}(144,44)(259,44){3}
//: {4}(260,44)(347,44)(347,36)(371,36){5}
//: {6}(372,36)(458,36)(458,36)(489,36){7}
//: {8}(490,36)(572,36){9}
input [3:0] A;    //: /sn:0 {0}(43,23)(173,23){1}
//: {2}(174,23)(288,23){3}
//: {4}(289,23)(404,23){5}
//: {6}(405,23)(521,23){7}
//: {8}(522,23)(565,23){9}
supply0 w10;    //: /sn:0 {0}(527,105)(591,105)(591,106)(601,106){1}
input Cin;    //: /sn:0 {0}(613,304)(464,304)(464,313){1}
//: {2}(462,315)(346,315)(346,318){3}
//: {4}(344,320)(235,320)(235,321)(225,321){5}
//: {6}(221,321)(104,321)(104,340){7}
//: {8}(106,342)(130,342){9}
//: {10}(102,342)(39,342)(39,133)(57,133)(57,143){11}
//: {12}(223,323)(223,338)(246,338){13}
//: {14}(346,322)(346,335)(368,335){15}
//: {16}(464,317)(464,335)(491,335){17}
output Cout;    //: /sn:0 {0}(1,165)(32,165)(32,166)(44,166){1}
supply1 w11;    //: /sn:0 {0}(612,232)(565,232)(565,231)(552,231){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(559,392)(512,392){1}
//: {2}(511,392)(390,392){3}
//: {4}(389,392)(267,392){5}
//: {6}(266,392)(152,392){7}
//: {8}(151,392)(60,392){9}
wire w6;    //: /sn:0 {0}(282,75)(282,69)(290,69)(290,61){1}
//: {2}(292,59)(304,59)(304,188)(282,188)(282,197){3}
//: {4}(290,57)(290,35)(289,35)(289,27){5}
wire w7;    //: /sn:0 /dp:1 {0}(230,253)(220,253){1}
wire w50;    //: /sn:0 {0}(391,348)(391,380)(390,380)(390,387){1}
wire w4;    //: /sn:0 {0}(133,139)(133,156)(73,156){1}
wire w25;    //: /sn:0 {0}(308,234)(324,234)(324,284)(379,284)(379,268){1}
wire w0;    //: /sn:0 {0}(194,105)(207,105)(207,166)(287,166)(287,144){1}
wire w22;    //: /sn:0 {0}(139,201)(139,187)(154,187)(154,60)(146,60){1}
//: {2}(144,58)(144,48){3}
//: {4}(144,62)(144,76){5}
wire w36;    //: /sn:0 {0}(528,193)(528,184)(542,184)(542,58)(525,58){1}
//: {2}(523,56)(523,35)(522,35)(522,27){3}
//: {4}(523,60)(523,67)(501,67)(501,72){5}
wire w20;    //: /sn:0 {0}(187,235)(200,235)(200,290)(244,290)(244,276){1}
wire w30;    //: /sn:0 {0}(428,230)(443,230)(443,291)(495,291)(495,273){1}
wire w37;    //: /sn:0 /dp:1 {0}(490,40)(490,46)(489,46)(489,56){1}
//: {2}(491,58)(512,58)(512,181)(500,181)(500,193){3}
//: {4}(489,60)(489,67)(467,67)(467,72){5}
wire w19;    //: /sn:0 {0}(510,142)(510,163)(429,163)(429,103)(419,103){1}
wire w23;    //: /sn:0 {0}(162,274)(162,316)(163,316)(163,326){1}
wire w54;    //: /sn:0 {0}(514,348)(514,380)(512,380)(512,387){1}
wire w21;    //: /sn:0 {0}(165,201)(165,185)(185,185)(185,62)(175,62){1}
//: {2}(173,60)(173,35)(174,35)(174,27){3}
//: {4}(173,64)(173,76){5}
wire w24;    //: /sn:0 {0}(153,355)(153,380)(152,380)(152,387){1}
wire w31;    //: /sn:0 {0}(403,197)(403,181)(422,181)(422,56)(407,56){1}
//: {2}(405,54)(405,27){3}
//: {4}(405,58)(405,66)(396,66)(396,73){5}
wire w1;    //: /sn:0 {0}(357,141)(357,302)(381,302)(381,319){1}
wire w32;    //: /sn:0 /dp:1 {0}(372,40)(372,56){1}
//: {2}(374,58)(387,58)(387,184)(371,184)(371,197){3}
//: {4}(372,60)(372,67)(363,67)(363,73){5}
wire w8;    //: /sn:0 {0}(259,144)(259,322){1}
wire w46;    //: /sn:0 {0}(269,351)(269,380)(267,380)(267,387){1}
wire w27;    //: /sn:0 {0}(252,197)(252,185)(271,185)(271,59)(262,59){1}
//: {2}(260,57)(260,48){3}
//: {4}(260,61)(260,69)(252,69)(252,75){5}
wire w28;    //: /sn:0 {0}(279,276)(279,322){1}
wire w33;    //: /sn:0 {0}(408,268)(408,309)(401,309)(401,319){1}
wire w41;    //: /sn:0 /dp:1 {0}(73,176)(87,176)(87,301)(134,301)(134,274){1}
wire w5;    //: /sn:0 {0}(305,107)(320,107)(320,165)(403,165)(403,141){1}
wire w38;    //: /sn:0 {0}(525,273)(525,309)(524,309)(524,319){1}
wire w9;    //: /sn:0 /dp:1 {0}(143,326)(143,311)(158,311)(158,139){1}
wire w51;    //: /sn:0 /dp:1 {0}(504,319)(504,311)(476,311)(476,142){1}
//: enddecls

  FA g4 (.B(w22), .A(w21), .Cin(w20), .Cout(w41), .S(w23));   //: @(120, 202) /sz:(66, 71) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Bo0<1 Bo1<0 ]
  mux g8 (.I0(w4), .I1(w41), .S(Cin), .Z(Cout));   //: @(57,166) /sn:0 /R:3 /w:[ 1 0 11 1 ] /ss:0 /do:0
  FA g3 (.B(w37), .A(w36), .Cin(w10), .Cout(w19), .S(w51));   //: @(447, 73) /sz:(79, 68) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Bo0<0 Bo1<1 ]
  //: joint g16 (w6) @(290, 59) /w:[ 2 4 -1 1 ]
  tran g26(.Z(w21), .I(A[3]));   //: @(174,21) /sn:0 /R:1 /w:[ 3 1 2 ] /ss:1
  //: joint g17 (w32) @(372, 58) /w:[ 2 1 -1 4 ]
  FA g2 (.B(w32), .A(w31), .Cin(w19), .Cout(w5), .S(w1));   //: @(340, 74) /sz:(79, 66) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>1 Bo0<1 Bo1<0 ]
  //: joint g23 (Cin) @(346, 320) /w:[ -1 3 4 14 ]
  //: input g30 (B) @(40,44) /sn:0 /w:[ 0 ]
  tran g39(.Z(w54), .I(S[0]));   //: @(512,390) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:0
  //: joint g24 (Cin) @(464, 315) /w:[ -1 1 2 16 ]
  FA g1 (.B(w27), .A(w6), .Cin(w5), .Cout(w0), .S(w8));   //: @(222, 76) /sz:(82, 67) /sn:0 /p:[ Ti0>5 Ti1>0 Ri0>0 Bo0<1 Bo1<0 ]
  tran g29(.Z(w36), .I(A[0]));   //: @(522,21) /sn:0 /R:1 /w:[ 3 7 8 ] /ss:1
  //: joint g18 (w31) @(405, 56) /w:[ 1 2 -1 4 ]
  mux g10 (.I0(w8), .I1(w28), .S(Cin), .Z(w46));   //: @(269,338) /sn:0 /w:[ 1 1 13 0 ] /ss:0 /do:0
  //: input g25 (A) @(41,23) /sn:0 /w:[ 0 ]
  FA g6 (.B(w32), .A(w31), .Cin(w30), .Cout(w25), .S(w33));   //: @(351, 198) /sz:(76, 69) /sn:0 /p:[ Ti0>3 Ti1>0 Ri0>0 Bo0<1 Bo1<0 ]
  //: input g35 (Cin) @(615,304) /sn:0 /R:2 /w:[ 0 ]
  FA g7 (.B(w37), .A(w36), .Cin(w11), .Cout(w30), .S(w38));   //: @(481, 194) /sz:(71, 78) /sn:0 /p:[ Ti0>3 Ti1>0 Ri0>1 Bo0<1 Bo1<0 ]
  mux g9 (.I0(w9), .I1(w23), .S(Cin), .Z(w24));   //: @(153,342) /sn:0 /w:[ 0 1 9 0 ] /ss:0 /do:0
  //: joint g22 (Cin) @(223, 321) /w:[ 5 -1 6 12 ]
  tran g31(.Z(w27), .I(B[2]));   //: @(260,42) /sn:0 /R:1 /w:[ 3 3 4 ] /ss:1
  //: supply0 g36 (w10) @(607,106) /sn:0 /R:1 /w:[ 1 ]
  tran g41(.Z(w46), .I(S[2]));   //: @(267,390) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:0
  tran g33(.Z(w32), .I(B[1]));   //: @(372,34) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g42(.Z(w24), .I(S[3]));   //: @(152,390) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:0
  tran g40(.Z(w50), .I(S[1]));   //: @(390,390) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:0
  mux g12 (.I0(w51), .I1(w38), .S(Cin), .Z(w54));   //: @(514,335) /sn:0 /w:[ 0 1 17 0 ] /ss:0 /do:0
  tran g28(.Z(w31), .I(A[1]));   //: @(405,21) /sn:0 /R:1 /w:[ 3 5 6 ] /ss:1
  tran g34(.Z(w37), .I(B[0]));   //: @(490,34) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  FA g5 (.B(w27), .A(w6), .new_port(w7), .new_port(w7), .Cin(w25), .Cout(w20), .S(w28));   //: @(231, 198) /sz:(77, 77) /sn:0 /p:[ Ti0>0 Ti1>3 Li0>0 Li1>1 Ri0>0 Bo0<1 Bo1<0 ]
  mux g11 (.I0(w1), .I1(w33), .S(Cin), .Z(w50));   //: @(391,335) /sn:0 /w:[ 1 1 15 0 ] /ss:0 /do:0
  //: joint g14 (w21) @(173, 62) /w:[ 1 2 -1 4 ]
  //: joint g21 (Cin) @(104, 342) /w:[ 8 7 10 -1 ]
  //: joint g19 (w37) @(489, 58) /w:[ 2 1 -1 4 ]
  //: joint g20 (w36) @(523, 58) /w:[ 1 2 -1 4 ]
  tran g32(.Z(w22), .I(B[3]));   //: @(144,42) /sn:0 /R:1 /w:[ 3 1 2 ] /ss:1
  //: supply1 g43 (w11) @(612,243) /sn:0 /R:3 /w:[ 0 ]
  //: output g38 (S) @(63,392) /sn:0 /R:2 /w:[ 9 ]
  FA g0 (.B(w22), .A(w21), .Cin(w0), .Cout(w4), .S(w9));   //: @(119, 77) /sz:(75, 61) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Bo0<0 Bo1<1 ]
  //: joint g15 (w27) @(260, 59) /w:[ 1 2 -1 4 ]
  tran g27(.Z(w6), .I(A[2]));   //: @(289,21) /sn:0 /R:1 /w:[ 5 3 4 ] /ss:1
  //: output g37 (Cout) @(4,165) /sn:0 /R:2 /w:[ 0 ]
  //: joint g13 (w22) @(144, 60) /w:[ 1 2 -1 4 ]

endmodule
