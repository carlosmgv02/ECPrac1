//: version "1.8.7"

module FullAdder2(A, Cin, B, Cout, S);
//: interface  /sz:(96, 63) /bd:[ Ti0>A(14/96) Ti1>B(51/96) Li0>Cin(26/63) Bo0<Cout(28/96) Bo1<S(61/96) ]
input B;    //: /sn:0 /dp:1 {0}(198,211)(186,211){1}
//: {2}(182,211)(159,211)(159,239){3}
//: {4}(157,241)(139,241){5}
//: {6}(159,243)(159,330)(199,330){7}
//: {8}(184,213)(184,305)(198,305){9}
input A;    //: /sn:0 {0}(136,206)(150,206){1}
//: {2}(154,206)(165,206){3}
//: {4}(169,206)(198,206){5}
//: {6}(167,208)(167,271)(198,271){7}
//: {8}(152,208)(152,300)(198,300){9}
input Cin;    //: /sn:0 {0}(143,304)(171,304){1}
//: {2}(173,302)(173,278){3}
//: {4}(175,276)(198,276){5}
//: {6}(173,274)(173,225)(281,225){7}
//: {8}(173,306)(173,335)(199,335){9}
output Cout;    //: /sn:0 {0}(412,321)(386,321){1}
output S;    //: /sn:0 /dp:1 {0}(302,223)(352,223){1}
wire w8;    //: /sn:0 {0}(219,274)(275,274)(275,287)(285,287){1}
wire w17;    //: /sn:0 {0}(306,290)(355,290)(355,318)(365,318){1}
wire w14;    //: /sn:0 {0}(220,333)(355,333)(355,323)(365,323){1}
wire w11;    //: /sn:0 {0}(219,303)(275,303)(275,292)(285,292){1}
wire w2;    //: /sn:0 {0}(219,209)(271,209)(271,220)(281,220){1}
//: enddecls

  //: input g8 (A) @(134,206) /sn:0 /w:[ 0 ]
  and g4 (.I0(B), .I1(Cin), .Z(w14));   //: @(210,333) /sn:0 /w:[ 7 9 0 ]
  //: joint g16 (A) @(152, 206) /w:[ 2 -1 1 8 ]
  and g3 (.I0(A), .I1(B), .Z(w11));   //: @(209,303) /sn:0 /w:[ 9 9 0 ]
  //: joint g17 (B) @(184, 211) /w:[ 1 -1 2 8 ]
  and g2 (.I0(A), .I1(Cin), .Z(w8));   //: @(209,274) /sn:0 /w:[ 7 5 0 ]
  xor g1 (.I0(w2), .I1(Cin), .Z(S));   //: @(292,223) /sn:0 /delay:" 2" /w:[ 1 7 0 ]
  //: input g10 (Cin) @(141,304) /sn:0 /w:[ 0 ]
  or g6 (.I0(w17), .I1(w14), .Z(Cout));   //: @(376,321) /sn:0 /w:[ 1 1 1 ]
  //: input g9 (B) @(137,241) /sn:0 /w:[ 5 ]
  //: joint g7 (A) @(167, 206) /w:[ 4 -1 3 6 ]
  //: output g12 (Cout) @(409,321) /sn:0 /w:[ 0 ]
  //: joint g14 (Cin) @(173, 276) /w:[ 4 6 -1 3 ]
  //: output g11 (S) @(349,223) /sn:0 /w:[ 1 ]
  or g5 (.I0(w8), .I1(w11), .Z(w17));   //: @(296,290) /sn:0 /w:[ 1 1 0 ]
  //: joint g15 (Cin) @(173, 304) /w:[ -1 2 1 8 ]
  xor g0 (.I0(A), .I1(B), .Z(w2));   //: @(209,209) /sn:0 /delay:" 2" /w:[ 5 0 0 ]
  //: joint g13 (B) @(159, 241) /w:[ -1 3 4 6 ]

endmodule

module FullAdder(A, Cin, B, S, Cout);
//: interface  /sz:(96, 73) /bd:[ Ti0>A(22/96) Ti1>B(63/96) Li0>Cin(30/73) Bo0<S(31/96) Bo1<Cout(61/96) ]
input B;    //: /sn:0 {0}(93,188)(27,188)(27,124){1}
//: {2}(29,122)(35,122){3}
//: {4}(25,122)(9,122)(9,125)(-12,125){5}
input A;    //: /sn:0 {0}(-12,110)(8,110)(8,117)(14,117){1}
//: {2}(18,117)(35,117){3}
//: {4}(16,119)(16,193)(93,193){5}
input Cin;    //: /sn:0 {0}(-13,143)(80,143){1}
//: {2}(82,141)(82,125)(91,125){3}
//: {4}(82,145)(82,163)(92,163){5}
output Cout;    //: /sn:0 {0}(165,179)(193,179){1}
output S;    //: /sn:0 {0}(112,123)(167,123){1}
wire w14;    //: /sn:0 {0}(56,120)(63,120){1}
//: {2}(67,120)(91,120){3}
//: {4}(65,122)(65,168)(92,168){5}
wire w2;    //: /sn:0 {0}(114,191)(134,191)(134,181)(144,181){1}
wire w5;    //: /sn:0 {0}(113,166)(134,166)(134,176)(144,176){1}
//: enddecls

  //: input g8 (A) @(-14,110) /sn:0 /w:[ 0 ]
  xor g4 (.I0(A), .I1(B), .Z(w14));   //: @(46,120) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  xor g3 (.I0(w14), .I1(Cin), .Z(S));   //: @(102,123) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  or g2 (.I0(w5), .I1(w2), .Z(Cout));   //: @(155,179) /sn:0 /w:[ 1 1 0 ]
  and g1 (.I0(Cin), .I1(w14), .Z(w5));   //: @(103,166) /sn:0 /delay:" 1" /w:[ 5 5 0 ]
  //: input g10 (Cin) @(-15,143) /sn:0 /w:[ 0 ]
  //: joint g6 (B) @(27, 122) /w:[ 2 -1 4 1 ]
  //: input g9 (B) @(-14,125) /sn:0 /w:[ 5 ]
  //: joint g7 (A) @(16, 117) /w:[ 2 -1 1 4 ]
  //: output g12 (S) @(164,123) /sn:0 /w:[ 1 ]
  //: joint g11 (Cin) @(82, 143) /w:[ -1 2 1 4 ]
  //: joint g5 (w14) @(65, 120) /w:[ 2 -1 1 4 ]
  and g0 (.I0(B), .I1(A), .Z(w2));   //: @(104,191) /sn:0 /w:[ 0 5 0 ]
  //: output g13 (Cout) @(190,179) /sn:0 /w:[ 1 ]

endmodule

module CPA(A, C4, B, Sout, C0);
//: interface  /sz:(140, 103) /bd:[ Ti0>B[3:0](86/140) Ti1>A[3:0](28/140) Li0>C0(46/103) Bo0<Sout[3:0](29/140) Bo1<C4(80/140) ]
input [3:0] B;    //: /sn:0 {0}(42,87)(158,87){1}
//: {2}(159,87)(332,87){3}
//: {4}(333,87)(511,87){5}
//: {6}(512,87)(675,87){7}
//: {8}(676,87)(737,87){9}
input C0;    //: /sn:0 {0}(37,243)(74,243){1}
input [3:0] A;    //: /sn:0 {0}(40,125)(102,125){1}
//: {2}(103,125)(282,125){3}
//: {4}(283,125)(455,125){5}
//: {6}(456,125)(542,125)(542,126)(627,126){7}
//: {8}(628,126)(738,126){9}
output [3:0] Sout;    //: /sn:0 {0}(15,461)(66,461){1}
output C4;    //: /sn:0 /dp:1 {0}(674,294)(674,366)(675,366)(675,376){1}
wire w6;    //: /sn:0 {0}(456,129)(456,200){1}
wire w7;    //: /sn:0 {0}(253,249)(243,249)(243,331)(155,331)(155,302){1}
wire w4;    //: /sn:0 {0}(115,302)(115,446)(72,446){1}
wire w0;    //: /sn:0 {0}(103,129)(103,202){1}
wire w3;    //: /sn:0 {0}(283,129)(283,137)(282,137)(282,204){1}
wire w12;    //: /sn:0 {0}(600,240)(569,240)(569,329)(509,329)(509,295){1}
wire w10;    //: /sn:0 {0}(628,130)(628,167)(627,167)(627,203){1}
wire w1;    //: /sn:0 {0}(159,91)(159,99)(157,99)(157,202){1}
wire w8;    //: /sn:0 {0}(512,91)(512,200){1}
wire w17;    //: /sn:0 {0}(425,239)(401,239)(401,331)(332,331)(332,299){1}
wire w14;    //: /sn:0 {0}(638,294)(638,476)(72,476){1}
wire w11;    //: /sn:0 {0}(676,91)(676,109)(677,109)(677,203){1}
wire w15;    //: /sn:0 {0}(72,466)(468,466)(468,295){1}
wire w5;    //: /sn:0 {0}(333,91)(333,108)(334,108)(334,204){1}
wire w9;    //: /sn:0 {0}(293,299)(293,456)(72,456){1}
//: enddecls

  //: input g4 (A) @(38,125) /sn:0 /w:[ 0 ]
  tran g8(.Z(w3), .I(A[1]));   //: @(283,123) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  FullAdder g3 (.A(w6), .B(w8), .Cin(w17), .S(w15), .Cout(w12));   //: @(426, 201) /sz:(132, 93) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>0 Bo0<1 Bo1<1 ]
  //: output g16 (C4) @(675,373) /sn:0 /R:3 /w:[ 1 ]
  FullAdder g2 (.A(w10), .B(w11), .Cin(w12), .S(w14), .Cout(C4));   //: @(601, 204) /sz:(116, 89) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>0 Bo0<0 Bo1<0 ]
  FullAdder g1 (.A(w3), .B(w5), .Cin(w7), .S(w9), .Cout(w17));   //: @(254, 205) /sz:(123, 93) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>0 Bo0<0 Bo1<1 ]
  tran g10(.Z(w6), .I(A[2]));   //: @(456,123) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g6(.Z(w0), .I(A[0]));   //: @(103,123) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g7(.Z(w1), .I(B[0]));   //: @(159,85) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g9(.Z(w5), .I(B[1]));   //: @(333,85) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g12(.Z(w10), .I(A[3]));   //: @(628,124) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: input g5 (B) @(40,87) /sn:0 /w:[ 0 ]
  tran g11(.Z(w8), .I(B[2]));   //: @(512,85) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: output g14 (Sout) @(18,461) /sn:0 /R:2 /w:[ 0 ]
  concat g20 (.I0(w4), .I1(w9), .I2(w15), .I3(w14), .Z(Sout));   //: @(67,461) /sn:0 /R:2 /w:[ 1 1 0 1 1 ] /dr:0
  FullAdder g0 (.A(w0), .B(w1), .Cin(C0), .S(w4), .Cout(w7));   //: @(75, 203) /sz:(126, 98) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Bo1<1 ]
  //: input g15 (C0) @(35,243) /sn:0 /w:[ 0 ]
  tran g13(.Z(w11), .I(B[3]));   //: @(676,85) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1

endmodule

module CPA2(A, Sout, C4, C0, B);
//: interface  /sz:(40, 40) /bd:[ ]
input [3:0] B;    //: /sn:0 {0}(39,98)(141,98){1}
//: {2}(142,98)(312,98){3}
//: {4}(313,98)(482,98){5}
//: {6}(483,98)(674,98){7}
//: {8}(675,98)(755,98){9}
input C0;    //: /sn:0 {0}(41,234)(75,234){1}
input [3:0] A;    //: /sn:0 {0}(50,70)(93,70){1}
//: {2}(94,70)(267,70){3}
//: {4}(268,70)(436,70){5}
//: {6}(437,70)(628,70){7}
//: {8}(629,70)(746,70){9}
output [3:0] Sout;    //: /sn:0 /dp:1 {0}(50,407)(104,407){1}
output C4;    //: /sn:0 /dp:1 {0}(646,295)(646,361){1}
wire w6;    //: /sn:0 {0}(268,196)(268,74){1}
wire w13;    //: /sn:0 {0}(496,295)(496,412)(110,412){1}
wire w16;    //: /sn:0 {0}(629,194)(629,74){1}
wire w4;    //: /sn:0 {0}(112,296)(112,336)(226,336)(226,237)(250,237){1}
wire w0;    //: /sn:0 {0}(142,191)(142,102){1}
wire w3;    //: /sn:0 {0}(155,296)(155,392)(110,392){1}
wire w12;    //: /sn:0 {0}(419,237)(395,237)(395,342)(285,342)(285,296){1}
wire w18;    //: /sn:0 {0}(687,295)(687,422)(110,422){1}
wire w10;    //: /sn:0 {0}(483,197)(483,102){1}
wire w1;    //: /sn:0 {0}(94,191)(94,74){1}
wire w8;    //: /sn:0 {0}(325,296)(325,402)(110,402){1}
wire w17;    //: /sn:0 {0}(611,235)(572,235)(572,341)(455,341)(455,295){1}
wire w11;    //: /sn:0 {0}(437,197)(437,74){1}
wire w15;    //: /sn:0 {0}(675,194)(675,102){1}
wire w5;    //: /sn:0 {0}(313,196)(313,102){1}
//: enddecls

  //: input g4 (A) @(48,70) /sn:0 /w:[ 0 ]
  tran g8(.Z(w0), .I(B[0]));   //: @(142,96) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  FullAdder2 g3 (.A(w16), .B(w15), .Cin(w17), .Cout(C4), .S(w18));   //: @(612, 195) /sz:(119, 99) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Bo0<0 Bo1<0 ]
  //: output g16 (Sout) @(53,407) /sn:0 /R:2 /w:[ 0 ]
  //: output g17 (C4) @(646,358) /sn:0 /R:3 /w:[ 1 ]
  FullAdder2 g2 (.A(w11), .B(w10), .Cin(w12), .Cout(w17), .S(w13));   //: @(420, 198) /sz:(120, 96) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Bo0<1 Bo1<0 ]
  FullAdder2 g1 (.A(w6), .B(w5), .Cin(w4), .Cout(w12), .S(w8));   //: @(251, 197) /sz:(117, 98) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Bo1<0 ]
  tran g10(.Z(w5), .I(B[1]));   //: @(313,96) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: input g6 (C0) @(39,234) /sn:0 /w:[ 0 ]
  tran g7(.Z(w1), .I(A[0]));   //: @(94,68) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g9(.Z(w6), .I(A[1]));   //: @(268,68) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g12(.Z(w10), .I(B[2]));   //: @(483,96) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g5 (B) @(37,98) /sn:0 /w:[ 0 ]
  tran g11(.Z(w11), .I(A[2]));   //: @(437,68) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g14(.Z(w15), .I(B[3]));   //: @(675,96) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  FullAdder2 g0 (.A(w1), .B(w0), .Cin(C0), .Cout(w4), .S(w3));   //: @(76, 192) /sz:(125, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Bo1<0 ]
  concat g15 (.I0(w3), .I1(w8), .I2(w13), .I3(w18), .Z(Sout));   //: @(105,407) /sn:0 /R:2 /w:[ 1 1 1 1 1 ] /dr:0
  tran g13(.Z(w16), .I(A[3]));   //: @(629,68) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1

endmodule

module main;    //: root_module
wire w16;    //: /sn:0 {0}(412,202)(412,184)(400,184){1}
wire w13;    //: /sn:0 {0}(336,203)(336,129)(303,129){1}
wire [3:0] w6;    //: /sn:0 {0}(938,252)(938,243)(932,243)(932,212){1}
wire w7;    //: /sn:0 /dp:1 {0}(473,412)(473,365){1}
wire w25;    //: /sn:0 {0}(947,206)(947,103)(904,103){1}
wire [3:0] w4;    //: /sn:0 /dp:1 {0}(479,260)(479,229)(427,229)(427,208){1}
wire w22;    //: /sn:0 {0}(927,206)(927,160)(905,160){1}
wire w3;    //: /sn:0 {0}(836,296)(867,296){1}
wire w0;    //: /sn:0 {0}(355,307)(392,307){1}
wire w20;    //: /sn:0 {0}(826,207)(826,189)(814,189){1}
wire w19;    //: /sn:0 {0}(846,207)(846,133)(813,133){1}
wire w18;    //: /sn:0 {0}(836,207)(836,161)(814,161){1}
wire w12;    //: /sn:0 {0}(422,202)(422,156)(400,156){1}
wire w23;    //: /sn:0 {0}(937,206)(937,132)(904,132){1}
wire [3:0] w10;    //: /sn:0 /dp:1 {0}(898,252)(898,247)(841,247)(841,213){1}
wire w24;    //: /sn:0 {0}(917,206)(917,188)(905,188){1}
wire w21;    //: /sn:0 {0}(856,207)(856,104)(813,104){1}
wire w8;    //: /sn:0 /dp:1 {0}(316,203)(316,185)(304,185){1}
wire w27;    //: /sn:0 /dp:1 {0}(941,393)(941,344){1}
wire w17;    //: /sn:0 {0}(442,202)(442,99)(399,99){1}
wire w14;    //: /sn:0 {0}(346,203)(346,100)(303,100){1}
wire [3:0] w2;    //: /sn:0 {0}(896,344)(896,386)(895,386)(895,393){1}
wire w11;    //: /sn:0 /dp:1 {0}(326,203)(326,157)(304,157){1}
wire w15;    //: /sn:0 {0}(432,202)(432,128)(399,128){1}
wire [3:0] w5;    //: /sn:0 {0}(421,260)(421,234)(331,234)(331,209){1}
wire [3:0] w26;    //: /sn:0 {0}(422,365)(422,414){1}
//: enddecls

  led g4 (.I(w7));   //: @(473,419) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: switch g8 (w11) @(287,157) /sn:0 /w:[ 1 ] /st:0
  //: switch g16 (w17) @(382,99) /sn:0 /w:[ 1 ] /st:0
  //: switch g3 (w0) @(338,307) /sn:0 /w:[ 0 ] /st:0
  //: switch g26 (w25) @(887,103) /sn:0 /w:[ 1 ] /st:0
  //: switch g17 (w16) @(383,184) /sn:0 /w:[ 1 ] /st:0
  //: switch g2 (w13) @(286,129) /sn:0 /w:[ 1 ] /st:0
  //: switch g23 (w22) @(888,160) /sn:0 /w:[ 1 ] /st:0
  //: switch g24 (w23) @(887,132) /sn:0 /w:[ 1 ] /st:0
  concat g1 (.I0(w8), .I1(w11), .I2(w13), .I3(w14), .Z(w5));   //: @(331,208) /sn:0 /R:3 /w:[ 0 0 0 0 1 ] /dr:0
  //: switch g18 (w18) @(797,161) /sn:0 /w:[ 1 ] /st:0
  led g10 (.I(w26));   //: @(422,421) /sn:0 /R:2 /w:[ 1 ] /type:1
  concat g25 (.I0(w24), .I1(w22), .I2(w23), .I3(w25), .Z(w6));   //: @(932,211) /sn:0 /R:3 /w:[ 0 0 0 0 1 ] /dr:0
  CPA2 g6 (.B(w6), .A(w10), .C0(w3), .C4(w27), .Sout(w2));   //: @(868, 253) /sz:(113, 90) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Bo1<0 ]
  //: switch g7 (w14) @(286,100) /sn:0 /w:[ 1 ] /st:0
  //: switch g9 (w3) @(819,296) /sn:0 /w:[ 0 ] /st:0
  //: switch g22 (w20) @(797,189) /sn:0 /w:[ 1 ] /st:0
  //: switch g12 (w8) @(287,185) /sn:0 /w:[ 1 ] /st:0
  led g11 (.I(w2));   //: @(895,400) /sn:0 /R:2 /w:[ 1 ] /type:1
  led g5 (.I(w27));   //: @(941,400) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: switch g14 (w15) @(382,128) /sn:0 /w:[ 1 ] /st:0
  //: switch g21 (w21) @(796,104) /sn:0 /w:[ 1 ] /st:0
  //: switch g19 (w19) @(796,133) /sn:0 /w:[ 1 ] /st:0
  concat g20 (.I0(w20), .I1(w18), .I2(w19), .I3(w21), .Z(w10));   //: @(841,212) /sn:0 /R:3 /w:[ 0 0 0 0 1 ] /dr:0
  concat g15 (.I0(w16), .I1(w12), .I2(w15), .I3(w17), .Z(w4));   //: @(427,207) /sn:0 /R:3 /w:[ 0 0 0 0 1 ] /dr:0
  CPA g0 (.B(w4), .A(w5), .C0(w0), .Sout(w26), .C4(w7));   //: @(393, 261) /sz:(140, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Bo1<1 ]
  //: switch g27 (w24) @(888,188) /sn:0 /w:[ 1 ] /st:0
  //: switch g13 (w12) @(383,156) /sn:0 /w:[ 1 ] /st:0

endmodule
