//: version "1.8.7"

module main;    //: root_module
wire cIN;    //: /sn:0 /dp:1 {0}(290,35)(303,35)(303,105){1}
wire w0;    //: /sn:0 {0}(430,204)(430,210)(408,210)(408,160)(369,160){1}
wire w1;    //: /sn:0 /dp:1 {0}(78,104)(78,128)(244,128){1}
wire w14;    //: /sn:0 {0}(369,131)(418,131)(418,114){1}
//: {2}(418,110)(418,105){3}
//: {4}(416,112)(406,112)(406,98)(418,98)(418,85){5}
wire w2;    //: /sn:0 /dp:1 {0}(51,172)(51,185)(122,185)(122,155)(244,155){1}
//: enddecls

  led g4 (.I(w0));   //: @(430,197) /sn:0 /w:[ 0 ] /type:0
  led g3 (.I(w14));   //: @(418,78) /sn:0 /w:[ 5 ] /type:2
  //: switch g2 (cIN) @(273,35) /sn:0 /w:[ 0 ] /st:0
  //: dip g1 (w2) @(51,162) /sn:0 /w:[ 0 ] /st:0
  FA g10 (.Cin(cIN), .B(w2), .A(w1), .Cout(w0), .S(w14));   //: @(245, 106) /sz:(123, 68) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Ro0<1 Ro1<0 ]
  //: joint g5 (w14) @(418, 112) /w:[ -1 2 4 1 ]
  //: dip g0 (w1) @(78,94) /sn:0 /w:[ 0 ] /st:0

endmodule

module FA(Cout, S, Cin, B, A);
//: interface  /sz:(40, 40) /bd:[ Ti0>Cin(19/40) Li0>B(29/40) Li1>A(13/40) Ro0<Cout(32/40) Ro1<S(15/40) ]
input B;    //: /sn:0 {0}(160,154)(128,154)(128,104)(115,104){1}
//: {2}(113,102)(113,91)(123,91){3}
//: {4}(111,104)(95,104){5}
input A;    //: /sn:0 {0}(97,85)(102,85){1}
//: {2}(106,85)(113,85)(113,86)(123,86){3}
//: {4}(104,87)(104,159)(160,159){5}
input Cin;    //: /sn:0 {0}(99,123)(154,123){1}
//: {2}(156,121)(156,100)(170,100){3}
//: {4}(156,125)(156,129)(160,129){5}
output Cout;    //: /sn:0 {0}(277,142)(233,142){1}
output S;    //: /sn:0 {0}(275,100)(201,100)(201,98)(191,98){1}
wire w13;    //: /sn:0 /dp:1 {0}(212,144)(191,144)(191,157)(181,157){1}
wire w7;    //: /sn:0 {0}(160,134)(149,134)(149,91){1}
//: {2}(151,89)(153,89)(153,95)(170,95){3}
//: {4}(147,89)(144,89){5}
wire w12;    //: /sn:0 /dp:1 {0}(212,139)(191,139)(191,132)(181,132){1}
//: enddecls

  //: output g4 (Cout) @(274,142) /sn:0 /w:[ 0 ]
  and g8 (.I0(B), .I1(A), .Z(w13));   //: @(171,157) /sn:0 /delay:" 3" /w:[ 0 5 1 ]
  //: output g3 (S) @(272,100) /sn:0 /w:[ 0 ]
  //: input g2 (Cin) @(97,123) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(93,104) /sn:0 /w:[ 5 ]
  //: joint g10 (Cin) @(156, 123) /w:[ -1 2 1 4 ]
  xor g6 (.I0(w7), .I1(Cin), .Z(S));   //: @(181,98) /sn:0 /delay:" 4" /w:[ 3 3 1 ]
  and g7 (.I0(Cin), .I1(w7), .Z(w12));   //: @(171,132) /sn:0 /delay:" 3" /w:[ 5 0 1 ]
  or g9 (.I0(w12), .I1(w13), .Z(Cout));   //: @(223,142) /sn:0 /delay:" 3" /w:[ 0 0 1 ]
  //: joint g12 (A) @(104, 85) /w:[ 2 -1 1 4 ]
  xor g5 (.I0(A), .I1(B), .Z(w7));   //: @(134,89) /sn:0 /delay:" 4" /w:[ 3 3 5 ]
  //: joint g11 (w7) @(149, 89) /w:[ 2 -1 4 1 ]
  //: input g0 (A) @(95,85) /sn:0 /w:[ 0 ]
  //: joint g13 (B) @(113, 104) /w:[ 1 2 4 -1 ]

endmodule
